��   "�A��*SYST�EM*��V9.4�0341 1/�17/2024 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG4��DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S?ETHOST��wNSS* 8��D�FACE_N�UM? $DBG�_LEVEL�O�M_NAM� !��* D �$PRIMAR_�IG !$ALT�ERN1�<WAIT_TIA ��� FT� @�� LOG_8	�C�MO>$DNL�D_FI:�SUBDIRCAP��Ό �8 . 4� H�ADDR�TYP�H NGcTH��4�z �+LS�&$�ROBOT2PE�ER2� MASKn4MRU~OMG�DEV��PIN�FO.  $�$$X4�RC�M+� E�$| ��QSIZ�X�� TATU�SWMAILSE�RV $PLA�N� <$LIN><$CLU����<$TO�P$C�C�&FR�&�JE�C�!�%ENB �� ALAR�!BF�TP�/3�V8 }S��$VAR79�M ON,6��,6A7PPL,6PA� -5�B +7POR��#_|12ALERT�&��2URL }>�3ATTAC��0�ERR_THRO��3US�9�!�8R0CqH- YDMAXN�S_�1�1AMOD�2AI� o 2A�� (1APWD � � LA �0�N�D)ATRYsFDE�LA�C2@�'`AERcSI�1A�'RO�ICLK�HMt0�'� �XML+ \3SGF�RM�3T� XOU̩3Z G_��COP c1V�3Q�'C�2-5R_AU�� � XR�N1oUPDXPC�OU�!SFO ?3 
$V~Wo��@YACC�H�QS�NAE$UMMY1z�W2?BGED79�DG$$C["D̻o PR
!-4�R�DM*	  �$DIS����S�MB�
 T &�	BCl@DCI2�AI&P6EXP9S�!�PAR�8`�RANe@  �7aCL� �<(C�0�SPT9M
U� PWR�eh�{f�SMo !l5��!�"%�7YD�P�% 0%vR�0z&uP� _DLV�$|e�aNo3 Bj�xX_Y`�#Z_I�NDE,C�pOFF,� ~UR�yD�bs��   t 9�!<pMON��s\ c�vHOU�#EyA��v��v��LOC�A� Y$N�0H�_HE��PI�"/  dA`AR�P�&�1F�W_�~ �I!F�p;FAp�D�01#�HO_� �R�2P\`�S�TEL	% P K � !�0WO�` 5�QE� LV{:�2H#ICE�����P��  ����1���
��
�&�pS$Q/��  Y5�$X'0 O�
���F�����Z������$.� 2l�#`���<������� l���!`8����ܒe�l�@��L�;�p�����"�"5�_�`l�ߋ��� į֯�����0�B��T�f�x��� _FL�TR  N�w� U����������nxl�2�p�SH^}`D 1l� P_�"ρ��N�=� r�5ϖ�YϺ�}��ϡ� �����8���\�߀� Cߤ�g�y��ߝ����� "���F�	��|�?�� c����������� B��f�)���M���q� ��������,��P t7I�m�� ����Lp 3�W�{����/�6/�PPP_�L�A1��x!�1.q"0?/�p%1|�/�255.�%Lx/�܉�o#2v/��.� �/�/�/�/�&3 �/�.e0?&?8?J?�&4f?�.�0�?�?�?�?�&5�?�.U@OO(O:O�&6VO�.�@|O�O`�O�O��aP(�1������ �Q� ./�N<FANUCy_�_�_ �Qh_�_�_�_o%o7o Po]ooo�o@o�o �o�o�o�o�o#�N��o���mX|
�ZDT Status�o|�����}iRConn�ect: irc��//alert �~-�?�Q�c��w���@����Ǐُ��y��P�R���"htt}p�172.2� �94.39:60�63/zdtdata/��H�Z�l�~� ������Ɵ؟����u�$$c962b3�7a-1ac0-�eb2a-f1c�7-8c6eb5�7dbcdb  ?(test�V���ppasswo�rdY���������A�WX�_Rܢaz"Π bt�jucQYT,$��)��NQ�T� ;�x�_�������ҿ�� ����,��P�7�IϠ��mϪϑ��ۧ��^%�������N?ot SenD�V~n?PDM_DQ	^+~N"SMB 
J]��#���Oz߯ߕ� �I߈}$t��{\�_CLNT �2^)��4ct ���[|��?��0�u� T�f�������������;�M�,�q�B.S�MTP_CTRL' ��8P%l��� At������g����?[|[�N��EPPK�2���h�b����;SdUST�OM Kݫ�%$^P %$:TTCPIPE�K���ctXVUZR� ELV$��~i  H!T	��T��rj3_�tpt�jrOP�!KCL_d�$%>��!CRT���/VR�!CO�NS/esib�_smon/!