��  ���A��*SYST�EM*��V9.4�0341 1/�17/2024 A   ������CCBD_�DATA_T � <$CO�MMENT �$IMCMF_�CF  NE�NDWTWCWFkDBWCd	FGW�TOOL_NUM�W w   qN�~ _FR�w �TRQ��GAIN�$T{DC�$CJI �� T�$DSR`��	I VP�AA�CTL_�TI�$MOV�E_L�WG@D�RARHY& {4/PARM9� �N PEQE} ��K�D&��3�K�K�D_M����3�h�+ �F�STd��|SU�  � L$L�IMIT� �$INSERT_�DIhx$�AM�_F Us"SRBPҎ)P�'|I3/dBNR x �_d�!B=�'TE0��$b�!ALr�"�AE�'FV��#T�9�v!A2U�(UNJ8V� TVh5Uq8�GRAPH�'RE�TRYS�<1�<2~WEC_DDE&x� �1�7A_PO�0��2AN� �5#��TWL�3ALLT�0�VV'@�!�$VCp27@�2�$�2Ar6@LhP�HD_RA�X`ED�sAheA�GO"�@�� I�DVA_SWG2�@��Ah�@5EhA� LE� �D�MC�ORWPH��!-ASDFW�FY_j"�CP�APz1QTN_S�#�CNGFh$M�IN�@�"?A_ML�_LM�VEL_�CNST�C$AUT_RVbUnPk@3_TL�0TH�1�T��1XSRUDAMP_��O|PS OLSTOP_THRE�1�TAV~Ub �P�D�SRAA�TM�Y��V��QATTOSC_GGDW�E*e#lR�FORCE_O�u MOF\eeI ��LSU�TJUT�fRO�T� C�1� CRE�W~#u �a�eCHG�ZQ�D�dDP@�cV��P��aR�1-AINISH�s�I�`_q�D�a^W�SoT@u|�WZPOCITYjmZP�CNm D�0�Dv Pdv��dZQ�P�V�t��#]#e/w/�/�/�'� �% (�$WOR� y2>�V  I��2U"�qST�P ����C1H�B�ry�RV~�����N�y�Fty�A	CTy�CWA����36��_M׊DCPdy�IV���V��ˇWQ���~��^Q��RTN|a��T�̇�a~�rALGO_Sxr�$P�1�t��R�EV_IT�1��MU�D�0CCI�!8RvȕXIŗGAM !f[AAS̖�_O@�NTR�vF�`�TuR�V%�CNPFv�6�?P�D�lDCNC�0M[ <��`O9�C%Hq�L�y�FG���\U�~�OVMI�Ql�,;���IOêD�AƦ�����JTH^QPqA�V�ݧPDA�p܃�%�DSPPCCN�MONLS
�D�T��1@�T�V�@j�KgPGRc���RG�1 ���d��R��O�t��%TʼO��Rp2����V�M�&�PDU~2CCNAGWA�g�1�TH�S?ǱAM�M0�S_ǖS0�VRS1}ɄŁ�M����82
�OVK�v��PG���U���±�VLx�;���TqCi��y�TRS?`V��MG�CCQ���T�H�s1R�INDE�mA�`TM3P�ft�C�Cߤt�RG]�USPF8w�Ժ���k@ߥ�TWD����f��SR����1D��˵���E�^PK�PPz��CAXCP_P�B1�l�.�3SRߣ3�DIQ�3��?PZh�U�&��RT�Y��LUFFIXE�CREG�Q+u�ㄬ�ߣF�q�P+CM<�r��CNFCf��SEN� R���V����RTV�TMU˵RG:�:�t���&:�DUE�3�TY�_�$0��S����PW��̂��IPI�:�APHf@����V�:�N��
� P1�M����� RC����>��W�P� H;�H�PYCIȫ��CHL�p�CK`V��c��q�VA��ΆPULIĆWATQ�I�I�I��HIPJ K�gS�IZ�SJ�DIAM��"�`����__���F��13;��=Oq�5�T#_jQ^0�! �E&PD]�MVR�OU2�PERI�O��F1� ��2D�G��T?�TU�_AD��甸ȅTڒ��K�KȅK�CqL���*aADJ���Q_U^B��AaPTp�bF%�2F#REP�H!�}H!Wuz+y)�D��*DL�W�$�*Mܠm��'0�)G��)�+ lB
9�'��)/3%:�)`N3D;8m3�'VL�* �3�:�)�3�;8�3�:N�+P_B���
�#�A�=��<�0�<OV3ER�D�2IB]PO'	Fq�TID0 TIe ��b"��FR�G�@d�rH!C5P�)MN1b��D2�NUF��KT#OOO��EAT�A�E1NG�X?QORܓ|BxAL{'wW��F��SU�e�6S1��AU�XBD0� 4?$IMCM�P�Ҁ��[� q�P!��`�P_7AXS�� �q�S� �` 	 h�PPEx`���T^c �S��S^ac=�h�W�D	hz`�� oX�AXI
P 
 �T���T��U�eA<�P�P xa'�~b	$Izh�`�f*��S�GRn�Hw $�AE_U�p&��d�B�a�@U�[���E֐�fswDO�N�a$FO��B�R_PKGry` � �bpxaSp�ar�a%r�`-t�pLp-p$��Sq~�$�VF/��_FILT�`��mqȅ�s���rׅlQ$DY�N�U$j }wG�w	�t��t׃	�QKa�`�
4�$ �  �����  � &� &�B@S�ION�?  Y5�� �a�COM ?.�&?� 2 �`� ^�p���������ʏ܏ � ��$�6�H�Z�l� ~�������Ɵ؟��� � �2�D�V�h�z��� ����¯ԯ���
�� .�@�R�d�v������� ��п�����4�?���`11 3M���9�4�j�1τǟ  �×�? ?�  �ū�A   �ŗ��ʯ�@@�˄����'�-�.�� B���-ژ�����q�Cяի�F�@ �ի�=���<�ի�Dz  �իϠ��o�-�Jі��`��W��h�{ύϟ� ���υ����߯���/� A�S�e�����߭߿� ����)���+�l�� ��k͟�k�������:��c�A���  @A���� ���aBHi��s�C��F�  �� 
��B�?� m�n��A�`u�>���;�k�D���d2����//*-	EB"2=/f/x/�/ �/�/�/�/�/�/?� ��)>��+O?�s� ��?��f�D��? �?O�?F���8G��?�9�dGP#��>���Ol�����8�E>L��?�A8�2�?�<#�
��p��O+B��*FS2������ECR� �E@���D�u_\ {� 0�]~O�B��E $�_o%ooIo[of� =�k�c��D �
�O�o��D�o�o��3It$ $�4&>��B
�oQwA��4Q�os/vD@+���̿u.�����u�q$敕�u(�4$��u��{;�{�.�>��H���q5��/�8M�Y;�K==�@W�CB (h�}�������ŏ׏�
���*��:� `�G�������{̟ß@՟���&�8�J�	� n�Y���}����ү� ����}_k�,�C�U� g�y���7oѿ�e ��	����?���c�u� ����KϽ����_�1� ����W߹��ρߓߴ� �%�7ϥ�[ϭ�ϑ� �ϵ�����������=� s����OI.�m� �������! 3%��_iN��� ������// S/8J\n��� ���?+?=?S?a? s?�?�?]߻?	��/�/ �/�/'O9O?]OoOT? �O�O�O�O�O�O�O_ #_5_G_Y_k_a?�_�_ �_�_�_��O�O�O1o _(_:_yo�o�o�/_ �o�_�_�_�-?$o c�_Fo�_���� so��)�;�M�_�q� Vhz���s�� ��
��.��R�d� v�eo��������Ǐ� ���<�'�`����o �_����̟ޟ�OA� &��+�=�O�a�s�_ ����;��?����� '�9�K�]�o�!��� #�5�G�Y�k�-Ϗ��� W�i�ׯ����{�1� ��U�g�y����ϯ��� ӿ����I������ C�U�g�y��������� ������	��-?$� cukߙ)������� ���� 2D Vhz����/ /)/7/I/_/m/O� ߏ����/?� 3?E?*/i?{?�?�?�? �?�?�?�?OO/O%/ 7/eOwO�O'?�O�ߕ? k?�?�?�?�?OO_a_ /��O�_qOaO�O�� oo'o�O�O0_�O�o �o�o�oI_�o�o�o #5G,o>oPoboto �oI��o�o�o�o�o �o(:L_pgy �����U��� 6�u�W��O~������� Əq?������I 7�I��?}��?��� ��������!�3�E� ��i�{ߩ���/�A� S�e�o�-�?�����џ �Q��Y�+�=�O�a� ���������߭���� �ߝ����+�=�O�}� s����������� ����9�K�A�o�T� f�x����������� ����,�>�P�b�t� ��u�����I�5 C%�ߵ^Ug� ��+	// ?/Q/ c/u/�/�/�/u�/�/ �/?���;?M?_?ُ �?=/k/��/�/�/�/ O%O7OIO�@?Od? [?m?g��O�O�O�?q? O�?W_i_{_�_#O�_ �_�_�_�_oo__ &_8_J_\_�_g_�_ �_�_�_�_�_o"o�? Fo=oOo|oso�o�o�o +��o�oK�-�?T fx��G/��ů ׯ鯿��A�S� g����e�����ӿ� ���ˏ-�/�Qς�� ���)�;�E��� ��������o�ݏ�� �%�7�}�[�m��q� �����Ϲ�������� �%�S��[�m�ߑ� �ߵߚ��������!� �E�*�<�N�`�r߱� ��ߺ��������� &�8�J�\�K������� ��������ߋo4� +�=�j������ ��'9K]o� f�������/ #/5/�Y/s�A�t W���/�/??Y� /U?:/1/O=�?�? �?�/G/�/k/-O?OQO cO�/�O�O�O�O�O�O �O�?�?�?O O�_�/ VO=OzOaO�O�O�O�O �O�O�/__%_R_I_ v_�_i_�_�_�_! oE*o<oNo`oroyc��$CCSCH_�GRP12 3�����a?&� �O�� ��a���ş韃> PqC�U�g�b��ݯ ����ӯ寸	��-� �o��&0��  �!������� ������h�F�X�j� ;�M��V�������.� ˿ݿ￵����7�I� O�m�ϑ��ϻ��� �����!�'�9�K�]� {ߊ��ߥϷ������� ���#�5�G�e�w�� ��������Ə�� ��C�:�s����ߩ� �������'9 K]o������ �����#5`�> _qT���� �V�/�I�/o �/��/��V�	? ?-???�c?u?�?�? �?�/�/�/�/�/?? �OA?(?:?w?^?�?�? �?�?�?�?��?+O"O 4OaOsO�O�_�O�O�O �O:/ _!o'_9_K_]_ o_F�(����������_ ��zo&o��:�L�^� 8o��ԟ����ʟܟ�o  ��$��_to�o�_�_ �_���Vohozo ��o�o�o�oz�o>� .@2��_Ə,�z� ��q���¯ԯ��
� ԟ.�@�%�d�v�\O�� ����п������� �!�3�r�C���{��� ����ÿտ����� \�n߀ߒߤ߆����� ���(�������j� |��Ϡ��6������� ��0�B�T�f�x��� ������������h� ,��5�t*�k�}� ����,����� �_�g�$� ,� //$/6/H/Z/ l/~/�/�/�/��� ����?/�'/M/ 4/q/X/�/�/�/��/ �/?�/
?7?I?[?�O ?j?�?�?�?�?�? O!O3O��_EO\n ����P��O�O~� �"�4�_X���|��� ����d_֏د��xOJ_ �O�Opo�O�_�o�o�o ,_>_P_�ot_�_�_�_ �_�_�_oo�VO ����b�G������� ���������(�:� L�>��g�����ʯ ܯ�ӟ���	�H�-� l�Q�c�u��������� ϯ��2�D�V�l�z� �Ϟϰ�vo��"?��¿ Կ�@�R�4�v߈�m� �߾���������*� <�N�`�r��zϨ�� ������
������J� �A�S�������.� �������FX=� |��_����� ��0BTfx� o������/� �#
G.k} �~������/ /1/�?U/@/y/�?�� ��/�/�/�/	?��ZO ??2oDoVohozo�o&� �?�?T�
�X?
,O. @Rdv�:O��� <?N?`?r?�?F_�?�O p_�_�?OO&O�_JO �OnO�O�O�O�_�O�O �O��bo��o8� \�n���������ȏڏ ����"��F�X�=� |����o��B�����͏ ߏ�0���'�9�K�]� o���������ɟ�� ,�B�P�b�x���h�/ �������ï�(�
� L�^�C��ϔϦϸ��� ���� ��$�6�H�>� P�~ߐߢ�@����o�� ��������)�h�z� H�Ư*����z߰ߚ/ �.�@��ߴ�I����� ������b���* <N`E�W�i�{��� ��b���������� ASe8��� ����n/+ O�/p�ߗ��� ���0?/__,_b� P_b_�ϖ/ �*��./ �/?oo(o:oLo^o �/�o�o�/$/6/H/Z/ l/~/�?FOXO�/�/�/ �/jO ?r?D?V?h?z? �O�?�?�?�o�o8_�o �o�_�_2DVh� ��������o �.�R�d�Z_��m ������� �!�3�E�W�i�{��� ���O���bo8�N� \�>��o�w�n����� ���D�"�4��X�j� |�������Ŀ����� �Ϯ��oT�f�x�� ��V���������ۿ� ,�>�P�bߜ�YϘ�}� tφπ�����ϊ� ߮�p����<��� ���� ��$�6��-� ?�Q�c�u�8���� ��������)�;�� _�V�h����������� D��%dF��m������$C�CSCH_GRP�13 3�����&� Ԕ_/�?�O�? 
OY.Oȿ����O �O�O��O"_�O__ *_�N_Pr_�U/ G]ku/3?E?f?� ��W?//1/C/�/ �?�?�/�/�/�_�_5O �O�_�_�Os?o"o4o ��XoC_|o�o�_�o�o �o\��o o0BYO flo~o�o�o��_� �o�o 2DVh z�����Ώ���� �(�?L�R�I�[��� ���ʟ5�� ���_ 6�H�Z�l�~������� Ưد���� �2�D� �Oh�z��O�������� گ�
��[�@ϛ�d� G�=���0�Z��ֿ�� ��񿛿-�N�`�r߄� 7Ϩߺ���������� �,�>�P�b����m� ߼ߣ��������(� :��C�p�g�y��� ����������E� fl�~��������OmO �/�/�/?/%?��Y k�O?�?�?}�?O �?�?O!O�EOGoiO ���+3AK	/ /</���-/�� �=�/as� wO��?q?�O�O�?�O __+_Y_O_Os_�_ jO�_�_����_�Oo 'o9o/?]oB_T_f_x_ �o�_�o�_�_�_�_o o,o>oPobo��� ���o���C�mo 1^U����� ��{�-�?�Q�c�u� ��������ϟ��؏ �)�;��?_�q�G�Y� z���o�����%� 7�q[���d�'�Q� ǿ���i�ǯq��E� W�i�{ύϟϱ����� ����޿���&�8� ��\�C�lϒ�y϶ϝ� ����������F�=� O�|ߎߠ���߯��� ��Y��0�B�T�f�x� ۏ�������� ���/�A��?U/g/y/ S��/�/�/�/�/�/�� ?_??������� �!��q����� ������Y 7I[M?���G/!� �?�/�?�?�?O/O%O �/IO[OmOO�O�/� �O�?�O�O_!_3_O *O<ONO�_rO�_�O�O �O�O�O�O__&_8_ wo�o�o�o�o�o�o�o �g��_oo+o� �yo���o��� '�9�K�]�o������� ��ɏ�o����#�5� O/�/�P���`����� ן���5os�1��� :�Q���������?��� G�]��-�?�џc�u� ��������Ͽ��Ưد ������2��V�h� O���s���¿Կß� ���%�R�d�v��� �υϾ���/�Y��� *�<�N�����w� ����k���/ O_��Oq�s��� �����?�ߓߥ� ���ߋ��������5� G�Y�k���������� ����/��1�#/5/ �Y/�}/b�/�/�/ �/?�/??1?C?U? g?/�?�?�/�?�?� �?�/�/ ??$?cOuO C?l?~?�?�?�?�?�? �?�?OM___q_�_�_ �_�_�_�OG�=��O�O �O_[omoO_�o�o�_ �o�o�o�o!3E Wi{��_�_�� ��o�%�o�o&	 J\n�����/_o ������a�s��� �����3���� ��9�K�]�o������� ��������ҟ䟧�� �,�>�%�b�I����� ��}�ίůׯ���(� :�L���p�[����ϵ� /�ܿ� ��$��ou� Z�M�_�q��O����A ��Eo%Os���G�I [m������ �i�{ύϟϱ����� �����/�A߯�e� �߉ߛ߭߿������ ��}�/A��8 w������� //+/=/"a/s/X �/�/���/���� �9?K?/B/T/f/x/ �/�/�/�/�/�/��5O GO)?�}O�O�O�? ��?�?�?�?1_C_�? g_y_^O�_�_�_�_�_ �_	o�O-o?oQoco�O /�o�o�o7��o�_�_ �?�_�_ o2oq�� ��?�o��o�o�oſ 7�I�[�!�od�o�� Ǐُ돁�!�3�E� W�i�{�`�r������� ��}�ޏŏ����8� �\�n���S������ ڟџ���"���F�1� j�������į֯������$CCSC�H_GRP14 �3���%��&� � ��S����=�Os� oȿڿ��������� �g�9�K�]�o�Bϓ� ���V�(Ϛό����� ��xߊ߫�
��.Ϝ� R�d�vψ�.� ����� ��������z��� %���Ugy??��� �����	�_? Ecu����� ��/)//AS ew������/ ??%?7?:/[?m?P� �?�/�/�/�/�/�?O z/3OEOG_"{O�O�O �O�O�O�O�O__/_ A_GOe_w_�_��_�_ ���O�O�O�O_1_Oo ao�O�o�/�o�_�_�_ u��o9?o6o�_ ro����|o�� �#�5�8M_q� ��I������ %��5�[�m��Ro�� ����������U�3� �W�B��o������ß ՟�������"�4� F�t�j�_����2��� ����¯�^�0�B�T� f������,���p� b�x�����N�`ρ�� ��r�(�:�L�^�� ���Ϧ���ʿ��
�P� ������:�L�^�p� ����^��������  �PO6�Zl~t� ������������  );M_q� ����
//./ R/d/*ψ/�dv� ��/?P*?<?�`? r?�?�?�?�?�?�?�? OO&O8O?\OnO�O �ߤO�O�?�?�?�O�? �?OF_X_j_|_��_ bOXO�Olo��o�O0o �O_�OH_�o�o�o�o �o�o�o,>#o 5oGoYoko}o@��o�o �o�o�o�o�o1C 2_^����� �L�	��-���_`� u��������� ?�Ϗ ���
��.�@��?t� ���ϬϾϘ���4� ��*�<��`�b��� �ԟ&�8���\�f�$� 6�W���ȟڟH���P� "�4�F�X���|����� ����ό�f/����� "�4�F�t�j�4ߎ�� ��������&?���0� B�T�f�x�]�o��� �������������#� 5�G�Y�k�}���� �(: �^� AL^p��� / /�6/H/Z/l/~/�/ �/�/�/�/�/�/? 2?D?V?h?z?��b/t/ �/�?�/�/�/O.O@O z�/vO8?.??�_�O �O�?_�?�?�?�_`_ r_�_O�_�_�_�_�_ oo�O__/_A_S_ w_^_�_�_�_�_�_ �_ooO)o4oFoXo jo�o�o�o"��o�o B�tO�?K]o�� >/����ί��� ��/J�\��ϔ���� ����ʿܿ� ��ď 6�8������П 2�<����z������� �ԏ&���
��.�t� R�d�v�h�z�쯞�0� �ϧ�����
��J�@� R�d�v߈ߚ߬�X��� �������<���3� E�W�iߨ��߱��� ��������/�A�S� ������������ ��o�o+�"�4�M�� �������0 BTfx���� �����//,/�P/ j�8kN��� �/?��P��L?// :/$�?�?�?H/>/�/ b/xO6OHOZO�/~O�O �O�O�O�O�O�?�?�? OO)O�_MO4OqO�O jO�O�O�O�O�O�/_ 
__5_@_m__�_�o �_�_�_�_t/!o3o EoWoio��o���� ����ڟ쟆 ��� j�o2�������į ֯�B��L�o�o �o�o�o�Џ�P bt����� ��J�(�:�L�>�P� t���@�}���ο� � ��(�:�L�^�p� ��g��ϸϝ������ ���	��-�?�~ߐ� aχϙϫϽ������� ��)��z��n�� ��������b�X_��� 
�7�v����߬����� ����*<N� r���8�t��� |o&��4�A$ ew����&�� "/�
o|/�/�/ f�8�/??0? �T?f?x?�?�?�?�? �/�/�/�/�/�/�O#? 
?G?.?@?}?d?�?�? �?��?�?�?OOCO UOgO�_�OvO�O�_�O�J�O	__-_?_HU��$CCSCH_G�RP15 3����jQ&� ���o^� 0������_��Roo @o�$�6�1oZ���~� �������o؟ڿ���_ mo�o�_�_�_�o�� �Ooaoso��o�o�o �ose�7�'9
� ���%�R�d�j���� �������͟��� <�N�`����������� ̿������,�J� Y�n�t���������ο ����4�F�X�j� |�Ϡ߲ߕ������ ���	�B�T��x�� ��g����������� ,�>�P�b�t������ ����a���/��.� @�#�d�v������ %��������OZ `~�{%��� �/�2/D/V/h/z/ }�������? /�	/F/-/j/Q/z/ �/�/�/��/�/�/? 0?B?T?�Ox?c?�?�? 	�?�O�?OO,O>O ���Ugy��O� I��O�Ow�	��-�_ Q���u�������]_Ϗ ѯ�qOC_�_�O�O�O �_�o�o�o%_7_I_�o m__�_�_Io�_�_ �_o�OO��I�[� @���������ٟ�� ����3�E�+?��{� `�����ï��̟ޟ ��A��e�J�\�n� ��������ȯگ�+� =�O�a�s�U��ϩ�oo ���������߿9�K� ��o߁�ϥ߷����� �����#�5�G�Y�k� }�bߡ����7����� �����C���:�L�� ��������������� ��?Q6�u��Q��� �����); M_q�hz�� ���/��� @'dv�w�a� ���//*/�?N/ 9/r/]/���/�/�/�/ �/?e�SO?+o=oOo aoso�o�?�?M��o �o�?'yK]o �3O����G?Ok? }??_�?�Oi_{_�_�? OO�_CO�OgOyO�O �O�_�O�O�O�%?[o �o��1�U�g�y��� ����yӏ���	�� k�Q�6�u������� ������Ə؏���;�  �2�D�V�h�z����� ����%�;�I�[� m��E_��������� ���!��E�W�<�{� �ϟϱ���������� �/�A�S�I�w߉ߛ� �߿��o�Ϲ������ �"�a�s�￯�ϻ� }�s������'��K� ��.�����������[� ����#5GY>� P�b�t�����[���� ��������:L^ M�ny�����  g/$H�/���� �������)?/ __%_7_I_[_�Ϗ/ �/#ٟ'/�_�/�_o !o3oEoWo	?{o}�/ ///A/S/Ow/�??O QO�/�/�/�/cO?k? =?O?a?s?�O�?�?�? �o�o1_�ou_�_+ =Oa����� ����o�'�K� ]�S_��x��� �������,�>� P�b�t�����ן��� ��1�G�U�7��� p�g�y������ٟ� -��Q�c�u������� ��Ͽ������ M�_�q���ϯ_}�S� ����Կ���7�I� ������Y�I��i�� ���σ�ߧϽ�{� ���1���������� �/��&�8�J�\�n� 1��y��������� �"�4��X�O�a�z� ��������=���� ]?��fx��� Y����?�?�?1�O 1O˿eϿ�_���w ��O�O�O	__-_� Q_c_��); MW/?'?���� 9?�A//%/7/I/�? m//�/�_�_O�_�_ �O�Ooo%o7oeo[o moo�o�o�o�o�_�o �o�_!3)OW<oNo `oro�o���o�o�o �o&8J\n ]?��я�1_��+� ��_��F�=�O�|��� ͟����'�9�K� ]�o�����]���ɯۯ �}��_#�5�G��k� %�S�y���i������� ��1�k�(�g�L�C� U�O�����ϫ�Y�� }�?�Q�c�u�ϙ߫� ��������������  �2�D��h�Oߌ�s� ���ߩ�����
�ݿ.� %�7�d�[���� �����3���<�N��`�r������$CC�SCH_GRP1�6 3������&� �cO��/u?�/�/ (�/��Rd�W?i? {?v�?�?�?�?�?�? �OoAO���$ ,:D//5/�� �&/�� ��/ |/Zl~OOaO?j? �O�O�?B/�O�O_� '_OK_]_cO�_�_�_ +��_�O�_�_o(?5o ;_M___q_�o�O�o�_ �_�_�_oo%o7oIo [oy�����o� ���!*WN ������Ϗџ�O� �)�;�M�_�q����� ����˟я����? 7�I�t?R�s���h��� ��ٯ�*��j3�� �]���)�����ÿɯ ��j����/�A�S�� wωϛϭϿ�¿׿� ����1���U�<�N� ��rϯϖϿ�����	� ܯ�?�6�H�u߇ߙ� ��ߨ�����N��5� ;�M�_�q��Z?<?� ��������(�:� �?N/`/r/L��/�/�/ �/�/�/��?_8?�� ���������� j�|���������� ���R0BTF? ���@/�?�?�/�?�? �?�?(OO�/BOTO9? xO�Op�ڏ�O�?�O�O _�,_O#O5OGO�_ WO�_�O�O�O�O�O�O �O__1_po�o�o�o �o�_�o�o�<_�_  o-o$o~��_�� Jo��� �2�D�V� h�z��������� ��
�|/.�@��(�I� ��>����П���� @o*���3���  {���8���@�ҟ�&� 8�J�\�n��������� ȿ����ѯ������ +��;�a�H���l��� ��Ϳ�������� K�]�o��ߓ�~ϷϢ� (������#�5�Gߪ ��Y�p����� d����/$6H"� l�����x�� �?/��^���߄��� �������@�R�d��� ����������(� �*�/jߠ�ov/ [�/�/�/�/�/�/� ?*?<?N?`?R��? {/�?�?�?�?O�/�/ ??\OA?�Oe?w?�? �?�?�?�?�?�?OF_ X_j_�_�_�_�_�_�� �_6��O�O�O�OTofo H_�o�o�_�o�o�o�o ,>Pbt� ��_����� �o�o^�/Ug�� ��ʏ_B ���	�  �Z�l�Q����s�� ,�������2�D�V� h�z������������� ˟ݟ����%�7�� [�B������������ Я���!�3�E���i� T�������(�տ��� ���on�S�F�X�j� |�����:����hO l�@�BTfx� �N���/P�b�tφ� ��Z���߄���� (�:ߨ�^߰߂ߔߦ� �������� ��v� (��L1p��� ���� //$/6/ �Z/l/Q�/�/���/ V����2?D?/ ;/M/_/q/�/�/�/�/ �/�/O.O@OVOdOvO �O�O|?���?�?�? �?*_<_O`_r_WO�_ �_�_�_�_�_oo&o 8oJo\oROdO�o�o�o T_�o���_�_�_�_o +o=o|�\�?>o� �o�o�o��0�B�T��o �o]�o���ҏ�v ��,�>�P�b�t�Y� k�}�������v�׏�� ����1��U�g�y� L��������ʟ��	� ���?�*�c������o ����ϯ��_D�)� �.�@�v?d�v�o�� o>�/B�����*� <�N�`�r�̿����ֿ 8�J�\�n�������Z� l�ڿ����~�4φ� X�j�|ώ��߲����� ����L������F Xj|����� ����0B'f xn������ //�#5GY k}�����?? �v�L?b?p?R/��� �/�/�/�/ OOX/6O HO-?lO~O�O�O�O�O �O�?�O_ _2_�?�� h_z_�_��_jO�O�/ �O�O�O_@oRodovo �/m_�o�_�_�_�� *�_�_3o�_�� ��Po����&� 8�J�/ASew� L�������� +�=�O�"os�j�|��� ��͏ߏ�X�� �9� x�Z��_��������ɟ�ҕ�$CCSCH�_GRP17 3������&� Ԩ� "��Ϻ���m�B��O ����ʯ�߮��߻��� 6���,�>��b�d ��%���i�[�q���� G�Y�z�ٯ���k�!� 3�E�W������ϟ��� ÿ���I߯������� ��$�6�H�/l�W�� ����������pO� 2DVm�z������ ��������"4 FXj|���� ��/	*/</�`/ f]o���/�/I ??O��J?\?n?�? �?�?�?�?�?�?�?O ?4OFOXO��|O�O�� �?�?�?�?�? O_0_ o?T_�x_[OQO�ODo n��_�Oo__�OA_ boto�o�oK_�o�o�o �ooo.o@oRodo vo��o�o�o�o�o�o �o*<N!_W� {����$��� &���_Y�z������� ��ȏ�߁�߿��� C�9��?m���ϥ� �ϑ���-����#�5� �Y�[�}���͟?�1� G�U�_��/�P����� ӟA���	��-�ӯQ� ��u�������ُυ� ������	��-�?�m� c�-߇��~߽��� ?���)�;�M�C�q� V�h�z���������� ����
��.�@�R�d� v��������! 3��W��3Eri ���/�//A/ S/e/w/�/�/�/�/�/ �/�/?�+?=?O?�� s?�?[/m/�/�?�/�/ �/O'O9OKO�oO1? '?x?;_e��O�?�O}? �?�?OY_k_}_�_�_ �_�_�_�_�_o�O_ _(_:_L_p_W_�_ �_�_�_�_�_ ooO �_-oZoQoco�o�o�o ��o�o�o�omO/D Vhz��ݏ��� ǯٯ�����/C�U� ��i�{���g����տ ���Ͻ�/�1�S�� ����ɟ+�5��� &��������͏�� ��'�m�K�]�o�a� ��[�5�Ϡ����� ��C�9��]�o߁� �ߥߗ��������� #�5�G�,�>�P�bߡ� ����߼�������� �(�:�L�������� ������	ϟ-{o� �-�?������� ��);M_q ��������/ /%/7/I/c�1Cd �/t���/�/?I� �E?/�N/eO�?�? �/�?S/�/[/qO/OAO SO�/wO�O�O�O�O�O �O�?�?�?�?O"O�_ FO-OjO|OcO�O�O�O �O�O�/�O__'_9_ f_x_�_�o�_�_�_ C?m/o,o>oPobo ��o��������ӟ� +��c�oc�� ��������ϯᯓ� ߕo�o�o�o�o�� �ɏۏI[m� ������C�!� 3�E�7�I���m����� v���ǿٿ���!� 3�E�W�i�{�'��ϱ� ������ݟߛ��� &�8�w߉�WπϒϤ� �����������"�a� s����������� [_Q_������o��� c������������ #5GYk}�� ��������9� ��:^p�� ����/��	 �_u/�/�/�1 G???)?�M?_?q? �?�?�?�?�/�/�/�/ �/�/�O??@?R?9? v?]?�?�?�?��?�? �?OO<ONO`O�_�O oO�O�_�OC�O__ &_8_���on_a�s��� �ߩ���U�_Y��9� �_o[o]�o������� ��o۟�o}_�_�_ �_�_�_�o��o1o CoUo�yo�o�o�o�o �o��o	���� C�U��L��������� ����	��-�?�Q� 6�u���l�������� Ưد����M�_�0� V�h�z�������¿Կ ����I�[�=ϻ��� �ߵߗ�1�'O������ �E�W��{��r߱� ������������A� S�e�w��C������� K_����������4� F������ϲ�� �������OK]o5 ��x����� #/5/G/Y/k/}/�/t ������?�� /�/L/3/p/�/�/ g�/�/�/�/�/?$? 6?�OZ?E?~?�O�?��?�?�?�?OE�$�CCSCH_GR�P18 3����9A&� ��g_-� Qc�O�!��O�O_ ��� _)�{�M�_� q���V_����ˏjO<_ �_�O�O�O�_�o�o�o _0_B_�of_x_�_�_ Bo4�_�_oُ� ��!�3�9��oi�{� ��Sϱ���՟��� �/���S�Y�w����� ���şן����(� =�C�U�g�y������� ��ӯ���'�9�K� N�oρ�do�ϫ����� �ؿ�#ߎ�G�Y�[� 6��ߡ߳��������� ��1�C�U�[�y�� ��0����������� ��3�E�c�u��ߙ��� ��������?)/� MS�J������� ���%7IL as����]/� ���9 Io ��f������ /#/i?G/2/k/V/�� �/�?�/�/�/�/?� �$o6oHoZo�?~o� �?�?F��o�o�o�?  rDVhz,O��� �@?O�Ov?�?�?�O b_t_�_�?OO�_<O NO`OrO_�O�_�O�O �O�?do�o�*� N�`�r�������r̏ ޏ����d�J�/� n������o�������� я��4��+�=�O� a�s������������ �0�B�$�f�x�>_�� Ɵx���������d� >�P�ԯtφϘϪϼ� ��������(�:�L� 1�p߂ߔ����ߠ� �������	��Z�l� ~��ʯ��v�l߽߀� �/ ��D��� ���\� ������������
 .@R7�I�[�m�� ��T���������� ��3EWF�0r� �����`/ A,��t���� �4�"?��O__0_ B_T_�ψ/�/�_�_ �_�/�_Hoo,o>oPo ?tov��o/�/:/L/ Op/z?8OJOkO�/�/ �/\O?d?6?H?Z?l? �O�?�?�?�o�*_�_ z� �_$6HZ� ~Ho������_ :� �D�V�h�z��� q�����
�� ��%�7�I�[�m�� ��П���
��*�<� N�Or��U�`�r��� ޯ�ҟ�&��J�\� n���������ȿڿ� ���"��F�X�j�|� �Ϩ_v������Ϲ�߿ �0�B�Tߎ�̿��L� BϓϪ��������� �Ϡ϶�t���*߼� ��������(��� 1�C�U�g�*��r�� �������	��-�� =�H�Z�l�~������� 6����V�߲�_ q���R����? �?�?OO*OĿ^p �_����O��O�O�O __&_�J_L�� �"�/FP/? ? ����2?�:// /0/B/�?f/x/�/|_ �_ O�_DO�_�O�_o o0o^oTofoxo�o�o �o�ol_�o�o�_, "OP�_GoYoko}o� ��o�o�o�o�o 1CUg����ʏ�� � ��$������?� 6�H�a���Ɵ����� � �2�D�V�h�z��� ����¯ԯ�܏�� .�@�ޟd�~OL�"�� b�����ǯ���_d� ȯ`�(��N�8���� ��\�R��v���J�\� n� ϒߤ߶������� ��������+�=� � a�H߅ߗ�~߻ߢ��� ���ֿ'��0�I�T� ���������, ���5�G�Y�k�}�(� ����/�/�/ ��/ ? ��4���O~��F� �?�?�?�?�?�?V O 2O`��������
 &��dv��/ ���^/< N`ROdO�/�O�OT? �?�O�O�O_4_*_<_ N_`_r_�_�_{O�_�_ �O�_o�/&o__/_ A_S_�o�ou_�_�_�_ �_�_�_oo+o=o,/ ���o O����o vOl�K���� �o��ҏ�����,� >�P�b�,��������� L��O�����:�� "�HU�8�y���ʯܯ � �:��6���$� �������z�(���L� � �2�D�گh�zό� �ϰ����Ϲ�˿ݿ� ����7��[�B�T� ��xϵ����Ϭ����� �3�*�W�i�{���� �������^���/��A�S�\��$CCS�CH_GRP19 3���~��&� �2?��rD/���� �f�!�3�T�&/8/J/ E�n/�/�/�/�/�/�� �/�O?��������� 	���c�u��� ����������yK );M?0?�9/f? x?~/�?�?�?�o�? �/O,O2?PObOtO�� �O�?�O�O�O�_
O O.O@O^_m?�_�O�O �O�O�O�O�O__*_ HoZolo~o�o�_�o�o ��o�_�_�_&ooV h�_����{?�� �
��.�@�R�d�v� �������Џ�u/� �C/!�B�T�7�x��� �����ޟ9o��ۏ ,�ί��n�t������� 9�˟����"�՟F� X�j�|���������ʯ ܯ� ���$���Z� A�~�e�����ƿؿ�� ����D�V�hϮ� ��wϰϛ�����
� �.�@�R�)//i{ �����]���	�/ /A�e��� ��q���?/��W� �������������� 9�K�]�������� ]���!���#�/c� �]/o/T�/�/�/ �/�/�/�?#?/G? Y??ϩ�?t/�?�?�? ��?�/�/??UO&? yO^?p?�?�?�?�?�? �?�? O?_Q_c_u_�_ iO�_�_���_O�O�O �O�OMo_o�O�o�o_ �o�o�o�o%7 I[m�vo�� �K���o�oW� N`����ÏՏ_ �����ş��e�J� ���e�������� �+�=�O�a�s����� |�������ğ֟���� �
�0��T�;�x��� ����u����ۯ�� ,�>���b�M���q��� ��ο����yog� (�?�Q�c�u�����3 ����a����; �_q��G߹�/ �[�-�ϑ�S�Ͽ� }����!�3ߡ�W� ��{ߍߟ߱������� ���9�o����_E* i{������ �////!oe/J �/�/�/�/�/��� �+?/O?4/F/X/j/ |/�/�/�/�/�/O'O 9OOO]OoO�O�OY�O ��?�?�?�?#_5_O Y_k_PO�_�_�_�_�_ �_�_oo1oCoUogo ]O�o�o�o�o�o���_ �_�_-�_$o6ou� ��?o��o�o�o� )�;� _��oB�o�� ��ˏݏo��%�7� I�[�m�R�d�v����� ��o�Џ�����*� �N�`�r�a������ ��ß���{�8�#� \�����o����ȯگ 쯗_=�"��'�9�K� ]�o�	o����7�/;� ����#�5�G�Y�k� Ϗ���1�C�U�g� )ߋ���S�e�ӿ��� 	�w�-��Q�c�uχ� �߫Ͻ�������E��� �� �?Qcu� �������� ); _qg�% ����//�
 .@Rdv�� ��/�/?%?3?E?[? i?K/�۟�/{/�/�/ �?O�//OAO&?eOwO �O�O�O�O�O�O�O_ _+_!?3?a_s_�_#O �_��OgO�O�O�O�O _Ko]o+�/_�om_ ]_�_}��o#�_�_ ,o�_����Eo� ����1�C�(: L^p�E���� �� ��$�6�H�o l�c�u�����Ə؏� Q����2�q�S��_z� ������mO����� ���E/3�E��Oy��O ����������� �/�Ae�w說� �+�=�O�a�k�)�;� ����ͯ߯M��U�'� 9�K�]��ρ������� �����������'� 9�K�y�o��������� ����������5G =�kP�b�t������ �������(: L^p�q���� E�/1/?/!�ﱏZ Qc��/�/'?? �;?M?_?q?�?�?�? q/�?�?�?O�/��7O IO[O՟O9?g?��? }?�?�?_!_3_E_ <O{_`OWOiOc��_�_ �_�OmO_�OSoeowo �o_�o�o�o�o�o �_o"o4oFoXo� |oco�o�o�o�o�o�o �OB9Kxo ���'����G� )��OP�b�t���������$CCSCH_�GRP1A 3����Á?&� �w�� ����ۿ�<�ϫ?f� x���k�}Ϗϊ���� ���������1�3�U� �Ɵ8�*�@�N�X�� (�I�����̟:��� �&�̯����n����� c�u��~ϫ߽���V� �����;�&�_�q� wߕ���??����� �%�<�I�O�a�s�� �������������� '�9�K�]�o���� ������/5 ,>kb��� ��/��/+/=/O/a/ s/�/�/�/�/�/�/� ??'?��K?]?��f/ �/�/|/�/�/�?�?>/ #O~GO*? ?q?_=� �O�?�O�?�?~?O1_ C_U_g_O�_�_�_�_ �_�O�O�O_!_3_E_ �oi_P_b_�_�_�_�_ �_�_oo�?&oSoJo \o�o�o�o��o�o�o �obO(I�Oas� �n�PϮ���ү�� ��/<�N���b�t��� `�����ο��϶� (�*�L����� �� $�.�����~����� �Ə؏����� �f� D�V�h�ZϨ�T��� �ϙ��������<�2� ��V�h�Mόߞ߄o� �߹���
���@�%� 7�I�[ߚ�k߾�ߵ� ���������!�3�E� �������������� ȟ&P���A�8�� �����^��" 4FXj|��� ����//��B/ T/*<]�/R�� �/�/??T�>? /� G/
O4�?�/�?L/�/ T/�/(O:OLO^OpO�O �O�O�O�O�O�?�?�? �?	OO�_?O&OOOuO \O�O�O�O�O�O�/�O �O)_ _2___q_�_�o �_�_�_�_<?�_o%o 7oIo[o��mo���� ����̟ޟx$�� 8�J�\�6��ү���� ȯگ��� �"��or �o�o���o�ԏ�� Tfx揜��� ��<��,�>�0�~o ��*���o�����ҿ ���ү,�>�P�b� t�f���Ϗ������� ������1�p�U� ��yϋϝϯ������� ��	��Z�l�~��� �������J_���� ���h�z�\������ ������
.@R dv������� �2� 3r Ci{����V /��4?n/�/e �/"�*@?�/?"? �F?X?j?|?�?�?�? �/�/�/�/�/�/�O? �/9?K?2?o?V?�?�? �?��?�?�?�?O5O GOYO�_}OhO�O�_/ <�O�O__1_���o g_Z�l�~�������N �_�_|�2߀_2�ToV� h�z�������boԟֿ d_v_�_�_�_n�_�o ��o*o<oNo�ro �o�o�o�o�o��o ����<�Ώ`�E� ���������ޯ�� �&�8�J���n���e� ������ڿj�ѯ��� �F�X�&�O�a�s��� ������Ϳ߿�0�B� T�j�xߊߠ߮ߐ�*O  O��������>�P�2� t��kߪ�������� ��(�:�L�^�p�f� xߦ�����h������ ��	���-�?�Q��� p���R���������O DVh����q / ����/./@/R/ d/v/�/m��� ��?��/!//E/ ,/i/{/�/`�/�/�/ �/�/??/?�OS?>? w?�O�?�?�?�?�? O��X_=O0BT�� x�$��O(�R��VO �O*_,�>�P�b�t��� �O�����OLO^OpO�O �O�O�_no�o�O __ $_�oH_�_l_~_�_�_ �o�_�_�_܏�`� $���Z�l�~����� ��Ɵ؟���� �� D�V�;�z�������� ����˟ݟ�.���%� 7�I�[�m�������� ǯ�o�*����`�v� ��f� ��/������տ �&�l�J�\�Aπߒ� �߶������߶��"� 4�F����|���O ��~߬�ҿ������ T�f�x���Ŀ������ ���?,>��� G������d�� (:L^CU gy��`/��� ��?Qc6� �~�����/ l?)//M/�?n/��/�/�/�/�/�%�$C�CSCH_GRP�1B 3����1&� Լ6O�_�o o 2o�?Vo�߫?�?�?�o �o�o�?�oJ.@ R%Ovx��9?O}O o?�?�?�O[_m_�_�? �?O_5OGOYOkO_ o�_�O�O�O��]o �o���_8�J�\� "���k�����ڏ� ����"�(�F�X�j��o ��������ʏ��� �$�6�H�Z�l�~��� ����ү������ >�P�3_t�z�q����� ����]��(�*�� ^�pςϔϦϸ����� �� ��$�*�H�Z�l� �o�ߢ��o�������� ��2�D��h�ï�� o�e߶�X��/����� "����U�v������� _��������0� B�T�f�x���,���� ��������>P b5�k����� �8/:%��m��/�����/�'C ??)?�O�_3o%_�� I_�Ϟ/�/�/�_�_�_ �/�_�_o!oT/Eo? iok��o,/�/P/b/t/ �/�?NO`O�?�/�/�? rO(?:?L?^?p?�O�O �?�?�?�o�oP_�_�o �o�_�O+=Oas ^o��o����_ Q�K�]�t_��� ��������� )�;�M�_�q������� şן����#�1�C� &Og�m�d�v�����Ͽ �L�	��-��oQ�c� �_��������ȟ�� ���;�M�_�q�K� ���_����ѿ����� %�7�I�[߶��b�X� ��K�u�߱���� ����i�{���R��� ��������5�5�G� Y�k�}������� ��������1�C�U�(� ^�������������+ 	��?]`�� �����D�/ /�?�O(_O��>O�� ����O�O�O��O �O__I:_/^_` �_!�EWi{�/ C?U?�/���/g?/ //A/S/e/�?�?�/�/ �/�_�_EO�O�_�_�O �? o2oDoVohoS_�o �o�O�o�o�o�O�_o F�@RiOv|o�o�o �o�o���o0 BTfx����̏ ޏ����&�8�?\� b�Y�k�����įڟA� ���"��_F�X��O|� ��������֯���� �0�B�T�f�@ϊ��O ����Ư������,� >�Pϫ�t�W�M���@� j�Ϧ��
�ϫ��� ^�p߂ߔ�Gϸ����� �� ��*�*�<�N�`� r���ߨߏ��߳��� ����&�8�J��S�� w������� ���� �4�RU�v|����������	E��/ �?O?�3?���� ��?�?�?��?�?�? O>/OSOUowO �:L^p�8/J/ ����\/$6 HZ�/�/����O �O:?�?�O�O�?x/_ '_9_K_]_HO�_�_�? �_�_�_w?�O_;�5o Go^?koq_�_�_�_�_ �o�o�_oo%o7oIo [omoo�o���� ���-�/Q�WN `����Ϗ6�� ��O;�M��?q����� ���˟ݟ���%� 7�I�[�5���?���� ����ߟ��!�3�E� �i�L�B��5�_�տ ������������S�e� wω�<��Ͽ������� ����1�C�U�g�	� �ϝτ��Ϩ������� �-�?��H�u�l�~� �߽���������)� G�J�k�q�������F������/? /�(/��}������/ �/�/���/�/�/ ?3� $?��H?J_l?���/� A�S�e�-?��� ���Q+=O �����z?�?// �/�?�?�/m
OO.O @ORO=?vO�O�/�O�O �Ol/�?�?0�*_<_S/ `_fOxO�O�O�O�_�_ �O�O__,_>_P_b_ t_�_�o�o�o�o�o "FLoCoUo�o yo���+o����? 0�B��/f�x�~���o ��ҏ�����,�>� P�*�t��/}������� ԏ���(�:��o^� A�7�t�*�T�ʯ��� ��럕���H�Z�l�~� 1�����ƿؿ��� �&�8�J�\��π��� y�����ڿ��ӿ�"� 4��=�j�a�sόϲ� ��
��������<�?߀`�f�xߊߜ߮���G ��������/��o ��r���w�� �����(�/�� =/?Oa/ ���$�6�H� Z�t�"4�������� F��� �2�D��� z�����o/�/$��/ �/�b�/?#?5?G? 2/k?}?��?�?�?a �/�/%�O1OHUO[? m??�?�?�O�O�?�? �?O!O3OEOWOiO{O �_�_�_�_�_�_oo ��;oA_8_J_w_n_� �o _�o�o�/%7 �[mso��_�� ���o�!�3�E�� i��r����� ����/��_S�6�,� i��I߿������� ����=�O�a�s�&��� ����ͯ߯�	�	�� -�?�Q��u���n��� ��ϯ��ȯ��)��� 2�_�V�h��������� ݿȿ��1�4�U�[� m�ϑϣ���H���� �߸������_| g�yߚ�l~��ߴ ������24? V�����+�=�O�i� �)���߻���;��� ��'�9����o�� ��dv��� W��//*/</'`/ r/��/�/�/V�� �?&?=J?P/b/t/ �/�/�?�?�/�/�/? ?(?:?L?^?p?�O�O �O�O�O�O�O_��0_ 6O-O?OlOcO�o�_O �_�_�_�o,o�Po boh_�o�O�o�o�o�o �_(:�^� go�o�o}o�o�o� � �$�OH�+!^� >ϴ�z؏��� 2�D�V�h�������� ԟ׏����"�4� F��j�|�c�����ğ ���������'�T� K�]�v�������ү�� ��&�)�J�P�b�t�������I�����ϭ� �����O�qo\�n� ��a�s����ϩ����� �����')/K� ��� �2�D�^��� �ߞϰ϶�0�����
� �.ߴ��d�v߈�Y k�t�����L�� �1Ug�� ���K���	/ /2�?/EWi{� �/�/����// //A/S/e/�?�?�?�? �?�?�?O��%O+?"? 4?a?X?�_�O
?�O�O �O�_!_��E_W_]O {_�?�_�_�_�_�O�_ oo/o	So~�\_}_ �_r_�_�_�o�o t?= ooSo	�3�� oo��o�oto�o'�9� K�]���������ɏ ��o���)�;�ݟ _�q�X���|������� ����o�I�@�R� k������ǟ��ן�� ��?�E�W�i�{�����J��ʿܿ��t��� �߲?��f_Q�c���V� h�z�u��������� ��˿�@�߯��� �'�9�S��ߒϓ� ����%�ۿ����#� �ߋ�Y�k�}�N�`�� i������A����� &�J\��� �@����o�'� 4:L^p��� ���� $6 HZx/�/�/�/�/�/ �/�/��? //)/V/ M/�O�?��?�?�?�� OO��:OLOR?pO{/ �O�O�O�O�?�O __ $_�_H_s�QOrO�OgO �O�O�_�_�_oi/2o __H_�o(��od_�o �_�_i__.@R ov�����o�_ �o�o0ҏTf M�q����� ��_�>�5�G�`��� ��ޟ����̏����4�:�L�^�p�����K ����ѯ��i����ϧ/ ��[OF�X�y�K�]�o� j��ߥ߷��������� �5�ԟ����
�� .�H���χ������� �Я������π� N�`�r�C�U���^ߋ� ���6�������	�� �?�Q���u�����5� �����O���)/� A�S�e�w������� ������+=O m������ ο/KBw? �/��/�/�/���/? ��/?A?G/e?p�?�? �?�?�/�?�?OO�O =Oh�F?g?y?\?�?�? �O�O�O_^'_
O O =O�_��_YO�_�O�O ^OtOo#o5oGo�Oko }o�o�o�o�_�O�_�_ oo%o�Io[oBoo fo�o�o�o�o�o�o�O 3*<U{�ӏ ������)�/� A�S�e�w�