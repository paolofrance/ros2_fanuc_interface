��  ��A��*SYST�EM*��V9.4�0341 1/�17/2024 A   ����DCSS_C�PC_T 4 �$COMMEN�T $EN�ABLE  �$MODJGRP�_NUMKL\�  $UFR�M\] _VTX �M �   $�Y�Z1K $Z�2�STOP_T�YPKDSBIO�IDXKENBL_CALMD��USE_PRED�IC? �ELAY�_TIMJSPEED_CTRLKOVR_LIM? *p D� �L�0�UT�OOi��O��4&S. ǰ 8J\TC �u
!���\�� jY0 � � �CHG�_SIZ�$A�P!�E�DIS"�]$!�C_+{#�s%O#J�p 	]$J d#� �&s"�"{#�)�$��'�_SEEX�PAN#N�iG�STAT/ D�FP_BASE_ $0K$4�!� .6_V7>H�73hJ- � q}�\AXS\3UP�LW�7����a7r � < w?�?�?��?�?�x//	7ELEM/ T �&B.2�NO�G]@%CNHA��DF#� $DAT�A)he0  �PJ�@ 2� 
&P5 �� 1U*n   �_VSiSZbRj0jR(��VyT(�R%S{TR/OBOT�X�SAR�o�U�V$CUR�_��RjSETU~4"	 $d �P_MGN�INP_ASSe#�P B!� `CiH�77`e��.fXc1�CONF�IG_CHK`E_�PO* }dSHRS�T�gM^#/eOTH�ERRBT�j_G]�R�dTv �ku�dVALD_7h�e�4hT1r
0R HLH8t� 0  lt<NerRFYhH~t�5"�1� ��W�_Ag$R��UPH/ (G%Q�Qt�Q3?wBOX/ 8�@F!�F!��G �r��zTUIR>i@  ,�F��pER%@2 �$�p l�_�Sf�A�ZN/O 0 IF(@L�p��Z_�0�_�08?wu0  @�QWy�v	*��~4�$$�CL`  �S��!���Q��Q�VERSION��  Yw5�$' 2 ?�Q  (��r���&@"�o�����������������Ԓd��Cz  2����C���n� ��������ȟݯ�� �"�4�F�H�j���� ��֯ǿ������� 0�B�T�f�hύϜ��� ��ҿ���ϐ��,�>� P��tωߘϪ�d��� ������(�:�`�^� p߅��߸������� ��$�6�H�Z�o�~� ������������  �2�D�j�Xz���� ��������. @Rdy���� ���	//*<N �b/��/����/ �??&/8/J/\/n/ �?�/�?�/�/�?�/O O%O4?F?X?j?lO�? �O�?�?�?�O�O_!_ 0OBOTOfOxO�O�_�_ �O�O�_�Ooo�_>_ P_b_t_/o�_�o�_�_ �o�_�o+:oLo^o �o�o�o�4�o�o�  �'�6HZl~ ������������ #�5�D�V�h���|��� ��ԏ���
��1� @�R�d�v��������� П�����-�?�N� `�r��������̯ޯ ���)�;�J�\�n� �����϶���ڿ�� �%�7�I�X�j�|ώ� �߲����������� 3�E�T�f�xߊߜ߮� ����������/�A� ��b�t���S����� ������=O^� p����������X��  $9KZl~ ��������  !/G/Y/hz�� �/��/��
/?./ C?U?d/v/�/�/�/�? �/�?�/?O*??OQO cOr?�?�?<O�O�?�O �?OO)_8OM___nO �O�O�O�O�_�O�_�O _%o4_Io[omo|_�_ �_�_�o�_�o�_oBo 3"Wixo�o�o�o �o�o��/�> S�e������w� �����Џ:�,�a��s�������̏ʏ܋��$DCSS_CS�C 2����Q  P ����<�ݏ`�#��� ��Y���}�ޯ���ů &�8���\����C��� g�ȿ��������"�� F�	�j�-ώϠ�c��� ���ϫ����0���T� f�)ߊ�M߮�q��ߕ� �����,���P��t� 7��[�m������盿GRP 2�� ����	ԟU�@� y�d������������� 	��?*cN� r������ M8q\�� ����/�/7/ "/[/F//j/�/�/�/ �/�/�/?�/?E?0? i?T?�?�?�?|?�?�? �?�?	O/OOSO>OwO �O�OfO�O�O�O�O_ �O_=_(_a_s_�_P_ �_�_�_�_�_�_o'o�oKo �_GSTA�T 2��'���< ��G�������?����k�?\��?�ǿ D��>�7�-��"���CD8��D4�'��:`<��f��;K
s��ᰅ� ���_%?�  �a?�`�4��Z�����e;���ڷ�?���p��K	ߌ����i@���Y�TDD1�=y=�.�����?~�z��K5�a��U��Rp)�J����.�2Dt����\?bR(bs�\��/=F��~?cj�>��� �L�?ӿe>D>��y��G<쾁~k?�" �F�I��cj�����?��`��7�?-���z�C�ODP<�{�o�o �k�u��>�P���2�|� ��h���ď҉�i�a�� ��y�0��(�J� x�^����������ʟ ܟ��,���\�n���z� ��~���گ��0�� D��L�2�D�f���z� ��ʿ��¿ ����� H�J����ϼ�v�����������;���?a%��e% �?W �>������u��՗�� L.�s���B�>�D;%��C�f��m��(ߖ?��ᴨ?{7�O�ar��<o��ow�k1�>�6�?l���<�
�lȆ�>�E���Կ��C���D$9��z���\>���|?sa��sм��)6�h�D<��2,�sN�>������s>����>�Hl?jt��<�1���?�w
�sQ����O���^DC�
C���y�<�^h?|b���*��w	�=sQ�>��Y�>�Վ> L$�?s� B��4�DAh�C� "�4�F�X��������� �$����Z�l��T� ���ߞ��������� ��J0R�fx ��B��
<�@ ,v�~���� ����/0//8/ f/L/^/�/�/�/�/�/ ��&?X?\?n?H? �?�?ߜ��T�f�x� �ߜ߮��������� �,�>�P�b�t���? �?�?�?x_�_�?�_�_ �_�_�_o��/2o4O :ohoNo`o�o�o�o�o �o�o�o6d �_���_���� �$�ohN�|F��� j�|���̏��ԏ�� ��8��0�R����,� �����
��.�@� �?8_J_�?OO&O8O JO\O�O�O�O�O�O�O �O�O�O_"_d�v��� "��&��J�\�6�H� �Ϥ�>�����Я��� �����L�2�T߂�h� �߸ߞ߰��� �z�0� B�t�N�x�R�d���� �������� ��� :�h�N�p��������� ���������^�� J�����V�Կ 濌�����¯ԯ��� F��.�@�R�d�v��� ������ $��/ �/��/�/�/�/.?@? ��(j?lr?�?�?�? �?�?�?�?OO&OTO :OLOnO�O?�O�O? �O_�O _J_\_R?�O �_�O~_�_�_�_�_o �_o:o o2opoVoho �o�o�Od_�o,_�o0 Bfx�p/�/( :L^p���� ��� //$/6/H/ Z/���ZL�^�T ����n���ʟܟv_�o ���<�"�4�V��� j�������¯�֯� 
�8���h�z������� ��������<�"�P� �X�>�P�rϠφϨ� �ϼ�������&�T� V� ϖ�ȿ�����߸� ������� ���0�~�T�f�x� ��������ҏ���8� J�\���������0 
fx�`ߢ�� ����� ( V<^�r��� N//H"/L/&/8/ �/�/���/��/�/ �/�/?<?"?D?r?X? j?�?�?�?�?�?��/ 2Od/OhOzOTO�O�O *����`�r���� ���������&�8� J�\�n������O�O�O �O�o�o�O�o�o�o�o �/�?>@_Ft Zl������ �(�� �B�p��o�� ���o���ԏ�0� &t�Z���R���v��� ��؟��������D� *�<�^�����8�ί �������:�L�B���$DCSS_JP�C 25bB�Q ( D?`��������P��ݿ ���������[�*� i�Nϣ�r��ϖ��Ϻ� ���3���i�8�J� \߱߀��ߤ������ ��A��"�w�F�X�j� ���������+��� O��0�r���f�x��� ��������9] ,�P�t��� ��#�1k: �^������ �1/ //$/y/H/�/ l/�/�/�/�/	?�/�/ ??? ?2?�?V?�?z? �?�?�?�?O�?�?:O _O.O@O�OdOvO�O�O �O_�O%_�OI__m_ <_N_�_r_�_�_�_�_��_��j�Ss�w�L �_Woo{o��dFo�o jo�o�o�o�o�o3 �oW{BTf� ������A�� e�,���P���t����� ����Ώ���O��s� :���^�����ߟ��� ʟ'�� ��[���H� ��l�ɯ�����د 5���Y� �g�D���h� z�������¿��C� 
�g�.ϋ�Rϯ�v��� �ϬϾ��-���Q�� u�<ߙ�`߽߄��ߨ� ������M��&�8� J��n�������� ��7���[�"��F�X� j�����������!�� Ei0�T�x �������S w>�b����/�(dMODE�L 25kx\��
 <�c(_  �|( �/i/{/�/�/�/�/�/ �/�/F??/?|?S?e? w?�?�?�?�?�?�?0O OO+O=OOOaO�_�O [/�O�O_�O�O>__ '_9_�_]_o_�_�_�_ �_�_�_�_:oo#opo GoYo�o}o�o�o�o�o �o�O�O�O�o~�o gy������ 2�	��-�?�Q�c��� ����揽�Ϗ��� �d�;�M���5Gu� ����o�ݟ���%� r�I�[���������� ǯٯ&����\�3�E� W�i�{���ڿ��ÿ� �������j��S�e� �ωϛ��Ͽ������ ��f�=�Oߜ�s߅� �ߩ߻�������P� '�9��!�3�E�s�� [�����(����^�5� G�Y�k�}��������� ����1C� gy������  �����?Q�u �������/ R/)/;/�/_/q/�/�/ �/�/?�/�/<??%? 7?�?1_?q?�?�? �?O�?�?JO!O3OEO �OiO{O�O�O�O�O�O �O�OF__/_|_S_e_ �_�_�_�_�?o�?�_ �_To+o=o�oaoso�o �o�o�o�o�o> '9K]o��� ������#��_ ��oK�]�ʏ���� � ׏�����1�~�U� g�����������ӟ� 2�	��h�?�Q�c�u� ����o�������ӯ@� �)�v�M�_�q����� ����˿ݿ*���%� r�I�[Ϩ�ϑ��ϵ� ����&�������	� 7�I߶�1ߟ߱����� ��4���j�A�S�e� w����������� ��+�=�O���s��� ��m�߭���,�� '9K]���� �����^5 G�k}���� /��H/����#/5/ �//�/�/�/�/�/ ? �/	?V?-???Q?�?u? �?�?�?�?
O�?�?O RO)O;O�O_OqO�OY/ k/}/�O�O�O__`_ 7_I_�_m__�_�_�_ �_o�_�_Jo!o3oEo Woio{o�o�o�o�o�o �o�o�OX�O!3	 w������� ��+�=���a�s��� ������͏ߏ�>���'�t�K�]�o����$�DCSS_PST�AT ����ՑQ  �  ��� � (�-��Q���v� t�֐�������������Օ��ׯ	�ƔSETU�P 	ՙB�������:�T�Ϭu��d���������I�ƔT?1SC 2
-�����Cz����);�CP R�D�DNtφ�@�� ���ϝ�����(�:� L�^�p߂ߔߦ߸��� ���� ��$�6�H�Z� l�~���������� ��� �2�D�V�h�z� ��������������
 .@Rdv��� `ϵ��Ϩ�� 3EWi{��� ����////A/ S/e/w/�/�/�/�/�/ �/�/??+?=?O?a? s?�?�?�?�?�?�?�? OO'O9OKO]OoO�O �O�O�O�O��O�O_ $5_G_Y_(_}_�_�_ �_�_�_�_�_oo1o CoUogoyo�o�o�o�o �o�o�o	-?Q cu������ ���)�;�M�_�q� ��������ˏݏ�� ��O7�I�[�n_��� ��r�ǟٟ����!� 3�E�W�i�{������� ïկ�����/�A� S�e�w���������ѿ �����+�=�O�a� sυϗϩϻ������� ��'�9�K�]�,��� �ߦ�t����ߪ���� #�5�G�Y�k�}��� ������������1� C�U�g�y��������� ������	-?Q cu������ �);M_q ��d߹����/ /%/�I/[/m//�/ �/�/�/�/�/�/?!? 3?E?W?i?{?�?�?�? �?�?�?�?OO/OAO SOeOwO�O�O�O�O�O �O�O__+_=_O_a_ s_�_�_�_�_�_�_� oo'o:/Ko]ooo>o �o�o�o�o�o�o�o #5GYk}�� �������1� C�U�g�y��������� ӏ���	��-�?�Q� c�u���������ϟ� ���)��_M�_�ro @�����v�˯ݯ�� �%�7�I�[�m���� ����ǿٿ����!� 3�E�W�i�{ύϟϱ� ����������/�A� S�e�w߉ߛ߭߿��� ������+�=�O�a�����$DCSS_�TCPMAP  ������Q @ Ġ�ĠĠĠ���ĠĠĠĠ	�Ġ
ĠĠĠ�ĠĠ9�  �ĠĠĠĠ*ĠĠĠġĠUĠĠĠĠUĠĠ Ġ!ĠU"Ġ#Ġ$Ġ%ĠU&Ġ'Ġ(Ġ)ĠU*Ġ+Ġ,Ġ-ĠU.Ġ/Ġ0Ġ1ĠU2Ġ3Ġ4Ġ5ĠU6Ġ7Ġ8Ġ9ĠU:Ġ;Ġ<Ġ=Ġ�>Ġ?Ġ@�UI�RO 2�������������  $6HZl~� ������á��7��[m� ������/!/ 3/E/W/i/{/�/�/ <�/�/�/??/?A? S?e?w?�?�?�?�?�? �?�?OO�/=O�/aO sO�O�O�O�O�O�O�O __'_9_K_]_o_�_��_�_0O�_{�UIZ�N 2��	 �����
oo.o4�o \ono�oCo�o�o�o�o �o�o�o4FX' |��c���� ��0�B��f�x�G� ������ҏ������ �>�P�b�%������� y�Ο��򟵟�(�:� 	�^�p���E�W���ʯ���� ���_��UF�RM R��� ���Y�k�}������� ſ׿�����1�C� U�g�yϋϝϯ����π����	��-�>�T��>�f�x�Sߜ߮߉� ���߿�����>�P� +�t��a������ �����(�?�Q�^�p� �������������  ��6H#l~Y �������  2I�Vh��y ����
/�./@/ /Q/v/�/c/�/�/�/ �/�/�/?*?AN?`? �/�?�?q?�?�?�?�? OO�?8OJO%OnO�O [O�O�O�O�O�O�O_ "_9?F_X_�Oi_�_�_ {_�_�_�_�_o�_0o BoofoxoSo�o�o�o �o�o�o1_P b��s��� ���(�:��^�p� K�������ʏ܏��� �$�;H�Z���~��� k���Ɵ�����ן � 2��V�h�C�y��������ԯ���
��4���$VALD_CP�C 2 ����@�Q  ���b�5� S A�R���f�@����ɿۿr�0���yd���Cz  � ��*�&��]�l�~��� �ϴ��������� � 2�D�V�k�zόϡ߰� ��������
��.�0� R�g�v߈߾߯���� ������*�<�N�c� u�����������x� ��&�8�M\�q�� ��L������� "HFXm��� �����0 BW/f{/���/� �/�/�///,/R/@? b/w?�/�/�/�?�/�? �???(?:?L?aOp? �O�?�?�O�?�O�O_ O$O6O�OJ_lO�_�O �O�O�_�O�_�__ _ 2_D_V_h_z_�o�_�_ �o�_�o�oo.o@o RoTvo��o�o�o� ��	�*<N` r������Ϗ�� ���&�8�J�\�q��� ������p�ڏ̟�� "�4�F�l�j�|���� ��ğٯ�����0� B�T�f�{��������� տ�����,�>�P� v�dφ��Ϫ���ο�� ���(�:�L�^�p� �ߔϩ߸�������� �'�6�H�Z� �n�� ������������#� 2�D�V�h�z���� ��������1@� R�d�v�x������� ��-<N` r������� /)/�J\n� �/��/���/��/ %?7?F/X/j/�/�/�/ �?@?�/�/�??!O3O B?T?f?x?�?�O�?�O �?�?�OO_/_A_PO bOtO�O�_�O�_�O�O �Oo_+o=oL_^_p_ �_�_�o�_�o�_�_ o'9KZolo~o$ ��o��o�o�o�  5�G�Vhz��� �׏����1�C� U�d�v���������ӟ ��*��
�?�Q�`� r���������ϯ�� ��&�;�M��n��� ������,�