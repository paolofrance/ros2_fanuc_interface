��   (�A��*SYST�EM*��V9.4�0341 1/�17/2024 A 	  ����PASSNA�ME_T   �0 $+ �$'WORD � ? LEVEL � $TI- OUTT4&F/�� $SE�TUPJPROG�RAMJINST�ALLJY  $CURR_OަUSER�NU�M�STSTOP�_TPCHG �V LOG_P NT��N�  6 C�OUNT_DOW�N�$ENB_�PCMPWD� �$DV_� IN�� $C� CR5E��A RM9� =T9DIAG9(|�LVCHK >FULLM/��YXT�CNTD��MENU�A�UTO+�FG_wDSP�RLS��U�BURYBA�N��GI�eE�NC/  ~CRYPTE�  �4��$$CL(   ���[!�� d �P V� IONX(�  Y5��$DCS_CO�D?���_%�  W�'_� �/�(WS  Z*�� \ ��&�A91�"[!�	 
 $��=  0b!9 7<B?X?f?|?�?�?�? �?�?�?�?OO0O>O�TO���#SUP� � :�?$?�#Fp�KWO�O'; \�Q�O_
�� �V�[t&��j
��.4hOp_��.W�,_�� �V�U�YqIL�UGH 1[)/ � �)�_ oo/oAoSoeowo�o �o�o�o�o�'�_�o #5GYk}�� ����o���1� C�U�g�y��������� ӏ��	��-�?�Q� c�u���������ϟ� ����)�;�M�_�q� ��������˯ݯ�� �%�7�I�[�m���� ����ǿٿ����!� 3�E�W�i�{ύϟϱ� ����������/�A� S�e�w߉ߛ߭߿��� ������+�=�O�a� s�����������  ��'�9�K�]�o��� ��������������� #5GYk}�� ������%