��  ��A��*SYST�EM*��V9.4�0341 1/�17/2024 A   ����DCSS_C�PC_T 4 �$COMMEN�T $EN�ABLE  �$MODJGRP�_NUMKL\�  $UFR�M\] _VTX �M �   $�Y�Z1K $Z�2�STOP_T�YPKDSBIO�IDXKENBL_CALMD��USE_PRED�IC? �ELAY�_TIMJSPEED_CTRLKOVR_LIM? *p D� �L�0�UT�OOi��O��4&S. ǰ 8J\TC �u
!���\�� jY0 � � �CHG�_SIZ�$A�P!�E�DIS"�]$!�C_+{#�s%O#J�p 	]$J d#� �&s"�"{#�)�$��'�_SEEX�PAN#N�iG�STAT/ D�FP_BASE_ $0K$4�!� .6_V7>H�73hJ- � q}�\AXS\3UP�LW�7����a7r � < w?�?�?��?�?�x//	7ELEM/ T �&B.2�NO�G]@%CNHA��DF#� $DAT�A)he0  �PJ�@ 2� 
&P5 �� 1U*n   �_VSiSZbRj0jR(��VyT(�R%S{TR/OBOT�X�SAR�o�U�V$CUR�_��RjSETU~4"	 $d �P_MGN�INP_ASSe#�P B!� `CiH�77`e��.fXc1�CONF�IG_CHK`E_�PO* }dSHRS�T�gM^#/eOTH�ERRBT�j_G]�R�dTv �ku�dVALD_7h�e�4hT1r
0R HLH8t� 0  lt<NerRFYhH~t�5"�1� ��W�_A�$R� �TPH/ (G%Q��Q�Q3?wBOX/ 8�@F!�F!��G �r��suUI}Ri@  ,��F�pER%@2 {$�p l�k_Sf�A�ZN/� 0 IF�(@�p��Z_�0�_p�0?wu0  @�Q�Wyv	*��~4�$�$CL`  ����!���Q��Q��VERSION��  �Y5�$' 2 �?�Q  ((�r���&@"�o�����������������Ԓd��Cz  2����C��� n���������ȟݯ� ��"�4�F�H�j�� ����֯ǿ������ �0�B�T�f�hύϜ� ����ҿ���ϐ��,� >�P��tωߘϪ�d� ��������(�:�`� ^�p߅��߸����� ����$�6�H�Z�o� ~������������  �2�D�j�Xz�� ���������� .@Rdy��� ����	//*< N�b/��/��� �/�??&/8/J/\/ n/�?�/�?�/�/�?�/ OO%O4?F?X?j?lO �?�O�?�?�?�O�O_ !_0OBOTOfOxO�O�_ �_�O�O�_�Ooo�_ >_P_b_t_/o�_�o�_ �_�o�_�o+:oLo ^o�o�o�o�4�o�o � �'�6HZl ~���������� ��#�5�D�V�h���|� ����ԏ���
�� 1�@�R�d�v������� ��П�����-�?� N�`�r��������̯ ޯ���)�;�J�\� n������϶���ڿ� ��%�7�I�X�j�|� �ϐ߲��������� ��3�E�T�f�xߊߜ� �߰���������/� A���b�t���S��� ��������=O ^�p����������X �� $9KZl ~������� � !/G/Y/hz� ��/��/��
/? ./C?U?d/v/�/�/�/ �?�/�?�/?O*??O QOcOr?�?�?<O�O�? �O�?OO)_8OM___ nO�O�O�O�O�_�O�_ �O_%o4_Io[omo|_ �_�_�_�o�_�o�_o Bo3"Wixo�o�o �o�o�o��/� >S�e������ w������Џ:�,� a�s�������̏ʏ܋��$DCSS_C?SC 2����Q  P����<�ݏ`�#� ����Y���}�ޯ��� ů&�8���\����C� ��g�ȿ��������"� �F�	�j�-ώϠ�c� �χ��ϫ����0��� T�f�)ߊ�M߮�q��� �������,���P�� t�7��[�m������~�GRP 2��' ����	ԟU� @�y�d����������� ��	��?*cN �r������ M8q\� �����/�/ 7/"/[/F//j/�/�/ �/�/�/�/?�/?E? 0?i?T?�?�?�?|?�? �?�?�?	O/OOSO>O wO�O�OfO�O�O�O�O _�O_=_(_a_s_�_ P_�_�_�_�_�_�_o�'ooKo �_GST�AT 2��'�ߜ< ��G��<����?��I��O�?\���?�� �F�>�6�-������CD?8�D4���:`�<�f��;K�s�ᰅ������%?�  �a?�`4��Z�����e�;��۷�j�?��p��K������i@��jd�T,�D�1=y=�C����8�?~�6�K5�a��W��?~��J�e��D2Dt���ھ�?b�R�bsjp=�F��?ckI>���}�L�?�u�D>�9y��G;W��}�?$n�F����ckK���v�?�`��6?-����z�C?��DPp�{�o �o�k�u��>�P���2� |���h���ď҉�i�a ����y�0��(� J�x�^���������� ʟܟ��,���\�n��� z���~���گ��0� �D��L�2�D�f��� z���ʿ��¿ ���� �H�J����ϼ�v�����Ϭ�����;���?a%��e%� ?W �>��澛�u������ L.�s���B�>�D;%��C�f��m�ʿ(�?����{7�O�a�r�<o��ow�k�1>�6�?l���<�
�l�߆>�E�������C���D$�9�y���\>���|?sa���sм�)6�h��D<�2,�sN��>������s>����>�Hl?jt�<�1����?w
�sQ�񾂜O����^DC�
C����y<�^h?|�b޾*��w�	=sQ�>���Y>�Վ> �L$?s� B���4DAh�C��"�4�F�X����� �����$����Z�l� �Tϖ��ߞ������� ����J0R� fx��B��
<� @,v�~�� ������/0/ /8/f/L/^/�/�/�/ �/�/��&?X?\? n?H?�?�?ߜ��T� f�xߊߜ߮������ ����,�>�P�b�t� ���?�?�?�?x_�_�? �_�_�_�_�_o��/ 2o4O:ohoNo`o�o�o �o�o�o�o�o 6d�_���_�� ���$�ohN�| F���j�|���̏��ԏ ����8��0�R��� �,������
�� .�@��?8_J_�?OO &O8OJO\O�O�O�O�O �O�O�O�O�O_"_d� v���"��&��J�\� 6�HϒϤ�>�����Я ��������L�2�T� ��hߊ߸ߞ߰��� � z�0�B�t�N�x�R�d� ����������� � ��:�h�N�p����� ������������� ^��J����� V�Կ濌�����¯ԯ ���F��.�@�R�d� v��������� $ ��/�/��/�/�/�/ .?@?��(j?lr?�? �?�?�?�?�?�?OO &OTO:OLOnO�O?�O �O?�O_�O _J_\_ R?�O�_�O~_�_�_�_ �_o�_o:o o2opo Voho�o�o�Od_�o,_ �o0Bfx�p/ �/(:L^p�� ����� //$/ 6/H/Z/���ZL� ^�T����n���ʟܟ v_�o���<�"�4� V���j�������¯� ֯�
�8���h�z��� ������������<� "�P��X�>�P�rϠ� �Ϩ��ϼ������� &�T�V� ϖ�ȿ���� �߸������ �����0�~�T� f�x���������ҏ� ��8�J�\��������� 0
fx�`� �������  (V<^�r� ��N//H"/L/ &/8/�/�/���/� �/�/�/�/?<?"?D? r?X?j?�?�?�?�?�? ��/2Od/OhOzOTO �O�O*����`�r�� ����������� &�8�J�\�n������O �O�O�O�o�o�O�o�o �o�o�/�?>@_ FtZl���� ���(�� �B�p� �o�����o���ԏ �0�&t�Z���R��� v�����؟������� �D�*�<�^�����8� ί ������:�L��B��$DCSS_�JPC 25bB��Q ( D?`��������P ��ݿ��������� [�*�i�Nϣ�r��ϖ� �Ϻ����3���i� 8�J�\߱߀��ߤ��� �����A��"�w�F� X�j��������� +���O��0�r���f� x�����������9 ],�P�t� ����#�1 k:�^���� ���1/ //$/y/ H/�/l/�/�/�/�/	? �/�/??? ?2?�?V? �?z?�?�?�?�?O�? �?:O_O.O@O�OdOvO �O�O�O_�O%_�OI_ _m_<_N_�_r_�_�_��_�_�_��j�Ss��w�L�_Woo{o��d Fo�ojo�o�o�o�o �o3�oW{BT f������� A��e�,���P���t� ��������Ώ���O� �s�:���^�����ߟ ���ʟ'�� ��[� ��H���l�ɯ���� �د5���Y� �g�D� ��h�z�������¿� �C�
�g�.ϋ�Rϯ� v��ϚϬϾ��-��� Q��u�<ߙ�`߽߄� �ߨ�������M�� &�8�J��n������ �����7���[�"�� F�X�j����������� !��Ei0�T �x������ �Sw>�b�����/�(dMO�DEL 25ksx��
 <�}c(  �|(�/i/{/�/�/�/ �/�/�/�/F??/?|? S?e?w?�?�?�?�?�? �?0OOO+O=OOOaO �_�O[/�O�O_�O�O >__'_9_�_]_o_�_ �_�_�_�_�_�_:oo #opoGoYo�o}o�o�o �o�o�o�O�O�O�o ~�ogy���� ��2�	��-�?�Q� c�������揽�Ϗ� ���d�;�M���5 Gu�����o�ݟ�� �%�r�I�[������ ����ǯٯ&����\� 3�E�W�i�{���ڿ�� ÿϫ������j�� S�eϲωϛ��Ͽ��� �����f�=�Oߜ� s߅��ߩ߻������ �P�'�9��!�3�E� s��[�����(���� ^�5�G�Y�k�}����� ��������1 C�gy���� �� �����?Q �u������ �/R/)/;/�/_/q/ �/�/�/�/?�/�/<? ?%?7?�?1_?q? �?�?�?O�?�?JO!O 3OEO�OiO{O�O�O�O �O�O�O�OF__/_|_ S_e_�_�_�_�_�?o �?�_�_To+o=o�oao so�o�o�o�o�o�o >'9K]o� �������� #��_��oK�]�ʏ�� �� �׏�����1� ~�U�g����������� ӟ�2�	��h�?�Q� c�u�����o������� ӯ@��)�v�M�_�q� ��������˿ݿ*�� �%�r�I�[Ϩ�ϑ� �ϵ�����&����� ��	�7�I߶�1ߟ߱� ������4���j�A� S�e�w�������� �����+�=�O��� s�����m�߭���, ��'9K]�� ������� ^5G�k}�� ��/��H/���� #/5/�//�/�/�/�/ �/ ?�/	?V?-???Q? �?u?�?�?�?�?
O�? �?ORO)O;O�O_OqO �OY/k/}/�O�O�O_ _`_7_I_�_m__�_ �_�_�_o�_�_Jo!o 3oEoWoio{o�o�o�o �o�o�o�o�OX�O! 3	w����� ����+�=���a� s���������͏ߏ� >��'�t�K�]�o�����$DCSS_P�STAT ����ՑQ?    ��� � (�-��4Q���v� t�֐@��������������Օ⯐�ׯ	�ƔSE�TUP 	ՙBȘ�����:�T� Ϭu�d���������I��ƔT1SC 2
4-�����Cz�����)��CP R�D�DNtφ� @�ϼ��ϝ����� (�:�L�^�p߂ߔߦ� �������� ��$�6� H�Z�l�~������ ������� �2�D�V� h�z������������� ��
.@Rdv ���`ϵ��Ϩ� �3EWi{� ������// //A/S/e/w/�/�/�/ �/�/�/�/??+?=? O?a?s?�?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O��O �O_$5_G_Y_(_}_ �_�_�_�_�_�_�_o o1oCoUogoyo�o�o �o�o�o�o�o	- ?Qcu���� �����)�;�M� _�q���������ˏݏ ����O7�I�[�n_ �����r�ǟٟ��� �!�3�E�W�i�{��� ����ïկ����� /�A�S�e�w������� ��ѿ�����+�=� O�a�sυϗϩϻ��� ������'�9�K�]� ,��ߓߦ�t����ߪ� ���#�5�G�Y�k�}� ������������� �1�C�U�g�y����� ����������	- ?Qcu���� ���);M _q��d߹�� ��//%/�I/[/m/ /�/�/�/�/�/�/�/ ?!?3?E?W?i?{?�? �?�?�?�?�?�?OO /OAOSOeOwO�O�O�O �O�O�O�O__+_=_ O_a_s_�_�_�_�_�_ �_�oo'o:/Ko]o oo>o�o�o�o�o�o�o �o#5GYk} �������� �1�C�U�g�y����� ����ӏ���	��-� ?�Q�c�u��������� ϟ����)��_M� _�ro@�����v�˯ݯ ���%�7�I�[�m� �������ǿٿ��� �!�3�E�W�i�{ύ� �ϱ����������� /�A�S�e�w߉ߛ߭� ����������+�=��O�aＨ�$DCS�S_TCPMAP  ������Q @ UĠĠĠĠ���ĠĠĠ�Ġ	Ġ
ĠĠ�ĠĠĠ9� � ĠĠĠ�ĠĠĠĠTġĠĠĠĠUĠĠĠ ĠU!Ġ"Ġ#Ġ$ĠU%Ġ&Ġ'Ġ(ĠU)Ġ*Ġ+Ġ,ĠU-Ġ.Ġ/Ġ0ĠU1Ġ2Ġ3Ġ4ĠU5Ġ6Ġ7Ġ8ĠU9Ġ:Ġ;Ġ<ĠU=Ġ>Ġ?Ġ@�UIRO 2����������� �� $6HZl ~�������á��7��[m ������� /!/3/E/W/i/{/�/ �/<�/�/�/?? /?A?S?e?w?�?�?�? �?�?�?�?OO�/=O �/aOsO�O�O�O�O�O �O�O__'_9_K_]_�o_�_�_�_0O�_{�U�IZN 2��	 �����
oo.o 4�o\ono�oCo�o�o �o�o�o�o�o4F X'|��c�� ����0�B��f� x�G�������ҏ���� ���>�P�b�%��� ����y�Ο��򟵟� (�:�	�^�p���E�W� ��ʯ��� ���_��UFRM R������Y�k�}��� ����ſ׿����� 1�C�U�g�yϋϝϯ� ��������	��-�>�T��>�f�x�Sߜ� �߉����߿����� >�P�+�t��a��� ���������(�?�Q� ^�p������������ �� ��6H#l ~Y������ � 2I�Vh� �y����
/� ./@//Q/v/�/c/�/ �/�/�/�/�/?*?A N?`?�/�?�?q?�?�? �?�?OO�?8OJO%O nO�O[O�O�O�O�O�O �O_"_9?F_X_�Oi_ �_�_{_�_�_�_�_o �_0oBoofoxoSo�o �o�o�o�o�o1_ Pb��s� �����(�:�� ^�p�K�������ʏ܏ ����$�;H�Z��� ~���k���Ɵ����� ן �2��V�h�C�y� ������ԯ���
���4��$VALD_�CPC 2 ����@�Q�  ��b�5�O  A�R���f�����ɿۿr�0����d���Cz  ���*�&��]�l� ~����ϴ�������� � �2�D�V�k�zό� �߰���������
�� .�0�R�g�v߈߾߯� ����������*�<� N�c�u��������� ��x���&�8�M\� q����L����� ��"HFXm� ������� 0BW/f{/�� �/��/�/�///,/ R/@?b/w?�/�/�/�? �/�?�???(?:?L? aOp?�O�?�?�O�?�O �O_O$O6O�OJ_lO �_�O�O�O�_�O�_�_ _ _2_D_V_h_z_�o �_�_�o�_�o�oo .o@oRoTvo��o�o �o���	�*< N`r������Ϗ �����&�8�J�\� q���������p�ڏ̟ ��"�4�F�l�j�|� �����ğٯ���� �0�B�T�f�{����� ����տ�����,� >�P�v�dφ��Ϫ��� ο�����(�:�L� ^�pυߔϩ߸����� ����'�6�H�Z� � n�ߥ���������� �#�2�D�V�h�z�� ����������� 1@�R�d�v�x��� ������-< N`r����� ��/)/�J\ n��/��/���/ ��/%?7?F/X/j/�/ �/�/�?@?�/�/�?? !O3OB?T?f?x?�?�O �?�O�?�?�OO_/_ A_PObOtO�O�_�O�_ �O�O�Oo_+o=oL_ ^_p_�_�_�o�_�o�_ �_o'9KZolo ~o$��o��o�o�o � 5�G�Vhz� ���׏���� 1�C�U�d�v������� ��ӟ��*��
�?� Q�`�r���������ϯ ����&�;�M�� n���������,�