��   "�A��*SYST�EM*��V9.4�0341 1/�17/2024 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG4��DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S?ETHOST��wNSS* 8��D�FACE_N�UM? $DBG�_LEVEL�O�M_NAM� !��* D �$PRIMAR_�IG !$ALT�ERN1�<WAIT_TIA ��� FT� @�� LOG_8	�C�MO>$DNL�D_FI:�SUBDIRCAP��Ό �8 . 4� H�ADDR�TYP�H NGcTH��4�z �+LS�&$�ROBOT2PE�ER2� MASKn4MRU~OMG�DEV��PIN�FO.  $�$$X4�RC�M+� E�$| ��QSIZ�X�� TATU�SWMAILSE�RV $PLA�N� <$LIN><$CLU����<$TO�P$C�C�&FR�&�JE�C�!�%ENB �� ALAR�!BF�TP�/3�V8 }S��$VAR79�M ON,6��,6A7PPL,6PA� -5�B +7POR��#_|12ALERT�&��2URL }>�3ATTAC��0�ERR_THRO��3US�9�!�8R0CqH- YDMAXN�S_�1�1AMOD�2AI� o 2A�� (1APWD � � LA �0�N�D)ATRYsFDE�LA�C2@�'`AERcSI�1A�'RO�ICLK�HMt0�'� �XML+ \3SGF�RM�3T� XOU̩3Z G_��COP c1V�3Q�'C�2-5R_AU�� � XR�N1oUPDXPC�OU�!SFO ?3 
$V~Wo��@YACC�H�QS�NAE$UMMY1z�W2?BGED79�DG$$C["D̻o PR
!-4�R�DM*	  �$DIS����S�MB�
 T &�	BCl@DCI2�AI&P6EXP9S�!�PAR�8`�RANe@  �7aCL� �<(C�0�SPT9M
U� PWR�ehx{f3co l5��!�"%�7Y�P��% 0%vR�0&uP� _DLV�|e�a	No3 BjxX�_Y`�#Z_IND9E,C�pOFF� ~UR�yD�bs�   t �!<pMON��s c�vHOU�#EyA�v�x�v��LOCA� �Y$N�0H_H-E��PI"/ w dA`ARP�&4�1F�W_~ �2I!F�p;FA�D�01#�HO_� �R�2yP\`�S�TEL	%G P K  !v�0WO�` �Q�E� LV{�2�H#ICE������P��  ��)�1���
��
&�p�S$Q/� ? Y5�$'0 VO�
���F�����Z������$� 2l��b��<��� ���� l���!8����ܒe�l���L��;�p�����"�5�_�`l�ߋ���į֯ �����0�B�T�f��x��� _FLTRs  N�w� ���������nx�l�2�p�SH}`DW 1l� P_�"ρ��N�=�r�5� ��YϺ�}��ϡ���� ��8���\�߀�Cߤ� g�y��ߝ�����"��� F�	��|�?��c��� ���������B�� f�)���M���q����� ����,��Pt 7I�m���� ��Lp3� W�{���/�|6/�PPP_L�A�1��x!1."q"0?/�p%1�/�255.�%x/�܉�o#2v/�.�  �/�/�/�/�&3�/�.@e0?&?8?J?�&4f?��.�0�?�?�?�?�&5 �?�.U@OO(O:O�&6VO�.�@|O�O�O�O،�aP(�1������ Q� ./�N<FANUCy_�_�_�Qh_��_�_�_o%o7o P o]ooo�o@o�o�o�o@�o�o�o#�N�o����mX|
ZD�T Status��o|����}�iRConnec�t: irc�/?/alert�~-� ?�Q�c��w�������PǏُ��y�P�R~���"http��172.2� 94�.39:6063�/zdtdata/��H�Z�l�~��������Ɵ؟����u$$�c962b37a�-1ac0-eb�2a-f1c7-�8c6eb57d�bcdb  (�test�V��p�password Y���������AఅWX�_RܢazΠ �bt�jucQYT,$ ��)��NQ�T�;�x� _�������ҿ����� �,��P�7�Iφ�m�h�ϑ��ۧ�^%��������Not� SenD�V~?PD�M_DQ	^+N"SMB 
J]�#����Oz߯ߕ� I߈}$t�{\��_CLNT 2*^)��4ct��� [|��?��0�u�T�f� �������������;�M�,�q�B.SMT�P_CTRL 	��8P%l���At�� ����g���?[|2[�N��EPK�2ԑ��h�b����;SdUSTOM' Kݫ%$^P� %$:TTCPIPE�K���ctVUZR�� ELV$��i  H!T	�T���rj3_tp�t�jrOP�!K�CL_d�$%��!CRT��/VR��!CONS�/esib_s'mon/!