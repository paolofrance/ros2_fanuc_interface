��  Ij�A��*SYST�EM*��V9.4�0341 1/�17/2024 A   ����SBR_T �  | 	$S�VMTR_ID � $ROBO�T9$GRP�_NUM<AXIaSQ6K 6NFF�3 _PARAM�F	$�  �,$MD SPD�_LIT4&2�*  � ���4�$$C�LASS  ����������� VERSION��  �Y5�$'  1 ~� T����
CRX-10�iA/L���  �biS1/6�000-B 40�A��
H1 D�SP1-S1��	P01.039�,  	� � ,  �P�P �� �����G��
�����
=�����o������ ��H�  ������ ����� w �����}�//1/~C/ ��g��/��5ҍ��!��2�� A� :?����'bD� ��/�/�/�/�/�/?i&8?J?\?��� \j?�?�?�?&��D0BTA2^�"j|��,�� ��>����O�O�O�OP(�r8��Vj/|/�/pF�/r_@�_�_�_?�_��)B �_�_ol?~?GoYokoH�?�?2�?T3^�)B"O4JBOTLF��FhOzL��	�:� 9�O�Hf� UBw�������xZE��Ox��*h��f5y,_>_P_ b_+�=�O�a��_����	�����ŏ׏2o�����1���o0��`0.3�e1QZ4^4�o0F� �<@Q AF �����<���~���{\D���J�&zh��@�@����[&\%�7�xI�[�������/��(v�w�p� ���,2��n� �1|B����	��v�?����va�s�����f 0- ����HϿ�<��F�0j�J|�5^5�������¿�TCʟܟ� �v��w[� ����������P% E�����?��(v" ������ү�߭߿��� ,���P��+�=J�s�����["�4)"�|�6^6FϠ������~���������hHw�����ϡ��������R$���b����(v�T�f�xߊ�S ew��߭�����P�+=O&8�?����Z�q(nn�'�	��a����//&/ 8/J/\/n/�/�/�/�/��/�/�/�/?"?2<� 2?V?h?z?�?�?�?�? �?�?�?
OC�~(O ����O�O�O�O�O �O�O__0_B_T_f_ x_�_�_�_�_�_�_@? oo,o>oPoboto�o �o�o�oOJO<O`O rO:L^p��� ���� ��$�6� H�Z�l�~����_��Ə ؏���� �2�D�V� h�z��o����0 ��
��.�@�R�d�v� ��������Я���� �*�<�N���r����� ����̿޿���&� 8ϴ���P�ʟܟ� ���������"�4�F� X�j�|ߎߠ߲����� �����h�0�B�T�f� x����������@� r�d�-��Ϛ�b�t��� ������������ (:L^p��� ���� $6 HZl~����� �4�F�X� /2/D/V/ h/z/�/�/�/�/�/�/ �/
??.?@?R?d?v? ��?�?�?�?�?�?O O*O<ONO`O��xO �//�O�O__&_ 8_J_\_n_�_�_�_�_ �_�_�_�_o"o4o�? Xojo|o�o�o�o�o�o �o�ohO�O�OU�O �O������� ��,�>�P�b�t��� ������Ώ��<o�� (�:�L�^�p������� ��ʟ&��\n� H�Z�l�~�������Ư د���� �2�D�V� h�z�������¿Կ� ��
��.�@�R�d�v� ��������,�>�� �*�<�N�`�r߄ߖ� �ߺ���������&� 8�J�\︿����� ���������"�4��� �ϴ�}����ϲ����� ����0BTf x������� d�>Pbt� ������N�/ 
/������p/�/�/�/ �/�/�/�/ ??$?6? H?Z?l?~?�?�?�?�? "�?�?O O2ODOVO hOzO�O�O�O,//�O B/T/f/._@_R_d_v_ �_�_�_�_�_�_�_o o*o<oNo`oro�o�? �o�o�o�o�o& 8J\�O�O�O� _ _����"�4�F� X�j�|�������ď֏ �����0��oB�f� x���������ҟ��� ��v?�2���� ������ί���� (�:�L�^�p������� ��ʿܿ�J��$�6� H�Z�l�~ϐϢϴ��� ��T�F���j�|���V� h�zߌߞ߰������� ��
��.�@�R�d�v� ������������ �*�<�N�`�r����� ����(�:�& 8J\n���� ����"4F X��j����� ��//0/B/��g/ Z/�������/�/�/�/ ??,?>?P?b?t?�? �?�?�?�?�?�?OO r:OLO^OpO�O�O�O �O�O�O�O _|/n/_ �/�/�/~_�_�_�_�_ �_�_�_o o2oDoVo hozo�o�o�o�o�o0O �o
.@Rdv ���_:_,_�P_ b_*�<�N�`�r����� ����̏ޏ����&� 8�J�\�n����o���� ȟڟ����"�4�F� X�j�������� � �����0�B�T�f� x���������ҿ��� ��,�>Ϛ�b�tφ� �Ϫϼ��������� (ߤ���@ߺ�̯ޯ�� �������� ��$�6� H�Z�l�~������ ������X� �2�D�V� h�z�����������0� b�T�xߊ�Rdv ������� *<N`r�� �����//&/ 8/J/\/n/�/�/���/ �/$6H?"?4?F? X?j?|?�?�?�?�?�? �?�?OO0OBOTOfO ��O�O�O�O�O�O�O __,_>_P_�/�/h_ �/�/?�_�_�_oo (o:oLo^opo�o�o�o �o�o�o�o $�O HZl~���� ���X_�_|_E��_ �_z�������ԏ� ��
��.�@�R�d�v� ��������П,�� �*�<�N�`�r����� �����߯үL�^�p� 8�J�\�n��������� ȿڿ����"�4�F� X�j�|ώ�ꟲ����� ������0�B�T�f� x���毐�
��.��� ��,�>�P�b�t�� ������������ (�:�L���p������� �������� $�� �ߤ�m���ߢ�� ��� 2DV hz������ �T�
/./@/R/d/v/ �/�/�/�/�/�/>? �/t��`?r?�?�? �?�?�?�?�?OO&O 8OJO\OnO�O�O�O�O /�O�O�O_"_4_F_ X_j_|_�_�_??�_ 2?D?V?o0oBoTofo xo�o�o�o�o�o�o�o ,>Pbt�O �������� (�:�L��_�_�_���_ oʏ܏� ��$�6� H�Z�l�~�������Ɵ ؟���� �|2�V� h�z�������¯ԯ� ��
�f�/�"������� ��������п���� �*�<�N�`�rτϖ� �Ϻ�����:���&� 8�J�\�n߀ߒߤ߶� ��D�6���Z�l�~�F� X�j�|�������� ������0�B�T�f� x��������������� ,>Pbt�� ��߽�*�� (:L^p��� ���� //$/6/ H/��Z/~/�/�/�/�/ �/�/�/? ?2?�W? J?����?�?�?�? �?
OO.O@OROdOvO �O�O�O�O�O�O�O_ b/*_<_N_`_r_�_�_ �_�_�_�_�_l?^?o �?�?�?no�o�o�o�o �o�o�o�o"4F Xj|���� _ ����0�B�T�f� x������_*oo�@o Ro�,�>�P�b�t��� ������Ο����� (�:�L�^�p������ ��ʯܯ� ��$�6� H�Z����r����� ؿ���� �2�D�V� h�zόϞϰ������� ��
��.ߊ�R�d�v� �ߚ߬߾�������� ��0謹��ο�� �����������&� 8�J�\�n��������� ������H�"4F Xj|���� � R�D�h�z�BTf x������� //,/>/P/b/t/�/ �/���/�/�/�/?? (?:?L?^?p?�?��? �?&8 OO$O6O HOZOlO~O�O�O�O�O �O�O�O_ _2_D_V_ �/z_�_�_�_�_�_�_ �_
oo.o@o�?�?Xo �?�?�?�o�o�o�o *<N`r�� �������p_ 8�J�\�n��������� ȏڏ�Hozolo5��o �oj�|�������ğ֟ �����0�B�T�f� x����������ү�� ��,�>�P�b�t��� �����Ͽ¿<�N�`� (�:�L�^�pςϔϦ� �������� ��$�6� H�Z�l�~�گ�ߴ��� ������� �2�D�V� h��ֿ�������� ��
��.�@�R�d�v� �������������� *<��`r�� �����p� ���]������ ����/"/4/F/ X/j/|/�/�/�/�/�/ �/D�/?0?B?T?f? x?�?�?�?�?�?.�? �?dv�PObOtO�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_�_ ?�_�_�_ oo$o6o HoZolo~o�oO�?�o "O4OFO 2DV hz������ �
��.�@�R�d��_ ��������Џ��� �*�<��o�o�o���o �o��̟ޟ���&� 8�J�\�n��������� ȯگ����l�"�F� X�j�|�������Ŀֿ ���V��ό����� xϊϜϮ��������� ��,�>�P�b�t߆� �ߪ߼���*����� (�:�L�^�p���� ��4�&���J�\�n�6� H�Z�l�~��������� ������ 2DV hz��߰��� �
.@Rd�� ��������/ /*/</N/`/r/�/�/ �/�/�/�/�/??&? 8?�J?n?�?�?�?�? �?�?�?�?O"O~GO :O����O�O�O�O �O�O__0_B_T_f_ x_�_�_�_�_�_�_�_ R?o,o>oPoboto�o �o�o�o�o�o\ONO�o rO�O�O^p��� ���� ��$�6� H�Z�l�~�������o ؏���� �2�D�V� h�z����o՟0 B
��.�@�R�d�v� ��������Я���� �*�<�N�`���r��� ����̿޿���&� 8�JϦ�o�b�ܟ� � ���������"�4�F� X�j�|ߎߠ߲����� ������z�B�T�f� x������������ ���v� ��ϬϾφ� ������������ (:L^p��� ���8� $6 HZl~���� B�4��X�j�2/D/V/ h/z/�/�/�/�/�/�/ �/
??.?@?R?d?v? �?��?�?�?�?�?O O*O<ONO`OrO��O �O//(/�O__&_ 8_J_\_n_�_�_�_�_ �_�_�_�_o"o4oFo �?jo|o�o�o�o�o�o �o�o0�O�OH �O�O�O����� ��,�>�P�b�t��� ������Ώ����`o (�:�L�^�p������� ��ʟܟ8j\%�� �Z�l�~�������Ư د���� �2�D�V� h�z��������¿� ��
��.�@�R�d�v� �Ϛ����ϲ�,�>�P� �*�<�N�`�r߄ߖ� �ߺ���������&� 8�J�\�n�ʿ���� ���������"�4�F� X�����p�������� ����0BTf x������� ,��Pbt� ������/`� ����M/�����/�/�/ �/�/�/�/ ??$?6? H?Z?l?~?�?�?�?�? �?4�?O O2ODOVO hOzO�O�O�O�O/�O �OT/f/x/@_R_d_v_ �_�_�_�_�_�_�_o o*o<oNo`oro�o�o �?�o�o�o�o& 8J\n��O�O� _$_6_��"�4�F� X�j�|�������ď֏ �����0�B�T��o x���������ҟ��� ��,����u�� �����ί���� (�:�L�^�p������� ��ʿܿ� �\��6� H�Z�l�~ϐϢϴ��� ����F���|����� h�zߌߞ߰������� ��
��.�@�R�d�v� ����������� �*�<�N�`�r����� ��$����:�L�^�& 8J\n���� ����"4F Xj|����� ��//0/B/T/�� �����/��
�/�/�/ ??,?>?P?b?t?�? �?�?�?�?�?�?OO (O�:O^OpO�O�O�O �O�O�O�O __n/7_ *_�/�/�/�_�_�_�_ �_�_�_o o2oDoVo hozo�o�o�o�o�o�o BO
.@Rdv �����L_>_� b_t_�_N�`�r����� ����̏ޏ����&� 8�J�\�n�������  ȟڟ����"�4�F� X�j�|��
��ů � 2�����0�B�T�f� x���������ҿ��� ��,�>�PϬ�bφ� �Ϫϼ��������� (�:ߖ�_�R�̯ޯ� �������� ��$�6� H�Z�l�~������ �������j�2�D�V� h�z������������� ��t�f��ߜ߮�v ������� *<N`r�� ���(��//&/ 8/J/\/n/�/�/�/  2$�/HZ"?4?F? X?j?|?�?�?�?�?�? �?�?OO0OBOTOfO xO��O�O�O�O�O�O�__,_>_P_b_�%��$SBR2 1��%�P T0? � ���/�'� �&#�UPl�_�_�_oo%o 7oIo[omoo�o�o�o�R��o�_�_' 9K]o���� ���o��o�o5�G� Y�k�}�������ŏ׏�����z���"�n�8�m���� ����ǟٟ����!� 3�E�(�:�L������� ïկ�����/�A� S�e�H�Z�l�~���ѿ �����+�=�O�a�sυϗ�z�~i_���� ����'�9�K�]�o� �ߓߥ߷����ظ��� 
��.�@�R�d�v�� �������������� *�<�N�`�r������� ��������&
� �\n����� ���"4FX <f������ �//0/B/T/f/x/ �/n�/�/�/�/�/? ?,?>?P?b?t?�?�? �?�?�/�?�?OO(O :OLO^OpO�O�O�O�O �O�O�O�?_$_6_H_ Z_l_~_�_�_�_�_�_ �_�_o o_DoVoho zo�o�o�o�o�o�o�o 
.@R6ov� �������� *�<�N�`�r���h�� ��̏ޏ����&�8� J�\�n����������� ڟ����"�4�F�X� j�|�������į֯�� ̟��0�B�T�f�x� ��������ҿ���� ��>�P�b�tφϘ� �ϼ���������(� :��^�p߂ߔߦ߸� ������ ��$�6�H� Z�l�Pߐ������� ����� �2�D�V�h� z��������������� 
.@Rdv� ������� *<N`r��� ����/�&/8/ J/\/n/�/�/�/�/�/ �/�/�/?"?4?/X? j?|?�?�?�?�?�?�? �?OO0OBOTO8?J? �O�O�O�O�O�O�O_ _,_>_P_b_t_�_jO |O�_�_�_�_oo(o :oLo^opo�o�o�o�o �_�o�o $6H Zl~����� ��o� �2�D�V�h� z�������ԏ��� 
�� �@�R�d�v��� ������П����� *�<�N�2�r������� ��̯ޯ���&�8� J�\�n���d�����ȿ ڿ����"�4�F�X� j�|ώϠϲϖ����� ����0�B�T�f�x� �ߜ߮���������� �,�>�P�b�t��� �������������� :�L�^�p��������� ������ $6� ,�l~����� �� 2DVh Lv������ 
//./@/R/d/v/�/ �/~�/�/�/�/?? *?<?N?`?r?�?�?�? �?�?�/�?OO&O8O JO\OnO�O�O�O�O�O �O�O�O�?"_4_F_X_ j_|_�_�_�_�_�_�_ �_oo0o_Tofoxo �o�o�o�o�o�o�o ,>PbFo�� �������(� :�L�^�p�����x�� ʏ܏� ��$�6�H� Z�l�~����������� ���� �2�D�V�h� z�������¯ԯ�ʟ ܟ�.�@�R�d�v��� ������п����� ��&�N�`�rτϖϨ� ����������&�8� J�.�n߀ߒߤ߶��� �������"�4�F�X� j�|�`ߠ�������� ����0�B�T�f�x� �������������� ,>Pbt�� ������( :L^p���� ��� //�6/H/ Z/l/~/�/�/�/�/�/ �/�/? ?2?D?(/h? z?�?�?�?�?�?�?�? 
OO.O@OROdOH?Z? �O�O�O�O�O�O__ *_<_N_`_r_�_�_zO �O�_�_�_oo&o8o Jo\ono�o�o�o�o�o �_�o�o"4FX j|������ ��o�0�B�T�f�x� ��������ҏ���� �,��P�b�t����� ����Ο�����(� :�L�^�B��������� ʯܯ� ��$�6�H� Z�l�~���t���ƿؿ ���� �2�D�V�h� zόϞϰ��Ϧ����� 
��.�@�R�d�v߈� �߬߾���������� *�<�N�`�r���� ������������
� J�\�n����������� ������"4F*� <�|������ �0BTfx \������/ /,/>/P/b/t/�/�/ �/��/�/�/??(? :?L?^?p?�?�?�?�? �?�?�/ OO$O6OHO ZOlO~O�O�O�O�O�O �O�O_�?2_D_V_h_ z_�_�_�_�_�_�_�_ 
oo.o@o$_dovo�o �o�o�o�o�o�o *<N`rVo�� ������&�8� J�\�n��������ȏ ڏ����"�4�F�X� j�|�������ğ���� ����0�B�T�f�x� ��������ү���ڟ �,�>�P�b�t����� ����ο����(� �6�^�pςϔϦϸ� ������ ��$�6�H� Z�>�~ߐߢߴ����� ����� �2�D�V�h� z��p߰��������� 
��.�@�R�d�v��� ������������ *<N`r��� ������&8 J\n����� ���/"/F/X/ j/|/�/�/�/�/�/�/ �/??0?B?T?8/x? �?�?�?�?�?�?�?O O,O>OPObOtOX?j? �O�O�O�O�O__(_ :_L_^_p_�_�_�_�O �O�_�_ oo$o6oHo Zolo~o�o�o�o�o�o �_�o 2DVh z������� 
��o.�@�R�d�v��� ������Џ���� *�<�N�