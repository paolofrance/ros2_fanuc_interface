��   -�A��*SYST�EM*��V9.4�0341 1/�17/2024 A   ����CELL_G�RP_T   �� $'FRA�ME $M�OUNT_LOC�CCF_METH�OD  $C�PY_SRC_I�DX_PLATF?RM_OFSCt�DIM_ $BA{SE{ FSETC���AUX_OR�DER   ��XYZ_MAgP �� ��LENGTH�T�TCH_GP_M�~ a AUTORA�IL_4�$$�CLASS  O�����D���DVERSIO�N  �Y5�8LOO�R G��DD<Z$?���q���M,  1 <DYX< [�����Cu��i�����iO/a/s/�A/�/�/�/$ ��/�/�/	;�$MN�U>A>"�  	 <i!/Q?�A? ?e?w?�?�?�?�?�? �?�?3OO+OMO{OaO �O�O�O�O�O�O�O_�/_�5NUM  %��	a��!2�TOOL%?\ !
;?/�_��_�_ �__�_%oo=o[oAo Souo�o�o�o�o�o�o �o)W=_��s���~VcS[
nY!