��  ��A��*SYST�EM*��V9.4�0341 1/�17/2024 A�  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ��4�ADV_I�N� 0  0KO�PEN� CRO �%$CLOS\� %EDI�BA �"IO_CNV�� l� RAC��LO�MOD_wTYP@FIR��HAL�#IN_;OU�FAC� g�INTERCEP:fB: SIZ@!�LRM_RECO�N"  � ALM��"=!  �&ON\�!� MDG/ �$DEBUG1PA2d43AO� �o"��!_IF�� � $ENA�BL@�#� P dj�#UU5K51MA�h� 2�
� OG�|f Z0CURR_�1:P $�3LIN@�1:�4$�$AUSO[4�� OD/2$SEV�_AND_NOA��2TP8"�6�4�5��APPINFOE=Q/  �L ��0�1EA H �GD9EQUI�P 38@NA�M/0�\B_OV�R�$VERS�I� �!PCOU�PLEm  	 �$�!PP�1CESI0�2�G101"P�0�B
 � $�SOFT�T_I�D�3OTAL_E%Q00�1�@N" �@U SPI
 �0^�E�X�3CRE ]Dn�BSIGz@�O|�K�@PK_FII0�	$THKY�RWPANE�D ~� DUMMY1d�yT!1�U4�Q  ��AR�1R� � $TITI1� ��0�Td�T!0��T�P�T5�V6�V7
�V8�V9�W �U�W@Q�U�W�Q�U�W1�WU1�W1g1g2b~�SBN_CF�![6@$L!J� �; K2A_CMNT��$FLAGS�]�CHE["$�b_OPTzB � �ELLSETUP�  `8@HO,h@I PR�1%�c#�	qREPRx�0D�+�@�+r{3uHM�I MN<% UTO�BZ U�0� D9DEVIC&�STI_@�� �@�r3�dpB�d�"VA�L3ISP_UN9I��p_DO�v7�yFR_FP�%�1�3��A`s�C_W�A�t\q�OFF_��@N�DEL1�L��0�q�1<��r?�q=�SS?��`2QRU1��#Z�;QTB1��b�MO� 1�E "REM1�����wREV�BILǇ��!XI� ��R 7 � OD�`끿$NO�`M@�������/�"���� �/��PD��d p E R�D_E〘�$F�SSB+6�`KBD�_SE�uAG� G
#Ba"_��2��� VQ�{5�`X��C�P`q	_8"�@2�r�$!�S�]D6 P�AQ�#�B;���_OK8a��0m P_C� ���`t�U pLACI��!q>���� �qC�OMM� # $D :�P�P=�ٙz_�R'@�BIGALLOW�� (K�2]BPVAR���!	Q�#�BL�@� � ,�K�qΤ�`S��@M�_O]����C?CFS_UTӀ@��"�AS�'-�[pX�w��b@ 40I'MCM0�3S�p��i�ʀi H�_D�<$���G��MA� hT�IMPEE_F�������� ���ǳD_�ӵ÷�DθF��4�_8H��@ T8@|��|�DI��@w�H�� =�PA�C$I?�W�M��F�d7 X8@GR�@�z�M��NFLI�<�ü@UIRE�y4<$2� SWIT~$p0k_N�`S02CF�0�M�,C@S��D��!�Ħ`-�<�J�`J�tV%�k E���.�p p(ڗELBOF� �IշI�p@p0���3�0��� F�2����BA��r�1J1,��z _T!��3p���g3p��rxPVCz� D��CLLB�`P=$�����F��G�� ��0WARNM�p��HK�`���`\ � COR-�r�FLTR��TRA�TI T? � $A�CC�qm�0r�r�$ORI�o&��ReT��Sl���HG�0I��T���A�I��T�t��� � &3�aa�N�HDR�2�2�2!J; HS'�!�3"� �$�5"�6"�7"�8"�9��
��
 /B� @0TRQB7�$�f���A�����_Ul�����O�c  <0�ϒϤ�E3�nB��LLECΒ!>"MULTI�4�"�2QK2M�CHILQD^�@!��O�@TM�w "W�STYI29r��=��)2���x��^�c# |�0 E6$�0�¦�`�L!�6uTO �E�	EXT����2�B2"��_��$�@�	N�p&��ak� %2k�p%qp�r���s�]�o&W���A���M���I )% ]T}R� ' L8@�{e#I r<�A��$JOBç���;IGi ( d��/ /)'r��#�a�Ǽ�@��_MOR��7) tT�FL1�:RsNGUQ��TBA�� P��&���*p1�(D�#@0��!�0;P�p 5�"�*$������qh`1w�rJw�_Rh���Cz<Jz�8�<J��D1�º9)���"'P���P_?pLҴ7+ \8@RORpHF�@��IT
�@NOM����,D3s:B!ڲ5UlPP�� �0�E,�P���0��PI��RA��ќѳC�[���
$T���MKD3$@T��pUp�L���+�AH�r��T1�JE5A����ÀQ�ƌQ�ƘQ�CYNT|����PDBGD��2�-^"ޠPU�$j�0�������AX)���4�TAI�sBUFp\�[YQ�. ���ljV�`PI��-�@P�WM�XM�Y\P�V�F�WSIMQST}O
�$KEE8cPA�є �BRR�C+R�� P��/�`��M�ARGA��2{�FA9C����LEW�1G!@�0��(�:����C�$c0W���@pJB���?qDEC�jL��ex����%1 �֐�CHN��MP��#$G�@7wt�_PCC�U�1_FPCEPTCbvv�S��tw�C���V{���q2��JR|��/�SEGFR�`�IO�!:@ST��L3INn��sPV����P]T2 ��rb����r��Ԡ�1�3` +�?��_�� 2p���`��)�j�y��aSIZ##���t�T��@�����RS��.#�s�Ӧypp�pL��
PAp$�gCRC��)�CC�р&��pN�bq��br|�MINz�bqz1`��4�D�iC��C��	ҕu`א�P��� ޘEVޖ�:�F��_�uF��N@ �<��a�ֱh�K�L��AS2
QVSCAuPA��rP���4C{ �SF0p4e����r �4P!Ҵ5��	��O�o �g�Ӡ�m��0�VP��b���Rs�6� �������e���R@HANC$cLGO�=��Q$蠳ND=���AR�N�8�qہ����̳ME`�Ҏ�Ͳ�PǸRA��̳AZ���
��EO��FCT�q�`pBBr�!S�`|0ADIm�Om���"��!��_�O�O �#s�G3�!9�'BMP�t��Y&COq��AES����n�W�_��BAS##XYOZWPR ����!:�	gAR_L~ ��_7( V�C��,����LBB'$g���!b�cv�pCEEVр�>FORCERQ��x`a'���_AVG���֫�MOMo0������S��TP�����А��i�=���F�d�A�YLOAD�$EAR/Љt�35B_X�pxc1"��QR_FD�_ 8 Tw`IQ $�3e Ed6:�C�:�[MS+`U{
$���p��)7d���9�eRHEVI��
�f�,1_IDX� $�倒�@�1���&�A��@�`R_9H�P��: �� 3���W!�f�_���; �]0��qpM<�q�@$PL�A��M��z�!���qF�������_CU�C�20��:��!PL߰���0T� �U5`M
�Um��<CTITA{
%_1�qTR �� �= PAEGED��� �PDT[R�EMd2`AUTH?_KEY  ) �bAD� @J NO���"Z_��mC>v�
��C߱FNO_HEADE�a�<� E�d�Pph�'��Ut�� M�V�e`�md?p�"P|��uCIRTR4p$4�N�L���C�@��RJ%�
��Q:�1�c@
B��:�OR!��9�O��M��qUN�_OðF�$SYAS1�5d�:�X����V�C�pe�DBPX�WO͐ A� $�SK�A�R*�DBT���TRLBv�A�C�p�D�u���DJ$�4� _���Qm$���y'PL!��bWA�"�� �cD`a�'8Q����2{ UMMY9���"10��PDBd�C+"�QPR6�
��DKо�D� m��1$;q�$��7�L8!E?�ci�@F7?$�/�PCAGV?$���PENE�@T�ڢHu?�2�!REC�ORP2IH ��@L�D$LK�E$3�R��;�p1���q�_D���PROS��T~�W���P0���TRIG )FP�AUS'C�tETU�RN'B�MRX�U2��9��0EW��>p?SIGNAL���R�$LAW��E��F{$PE�G$P8�2�AH�@��PC�DSi�DOIи��2�1c���6GO_AWAY�BMO�q�����!C�S��CSCBۡJC �/q��G��`I�@@� �R7p��'��6S�R@\``ARGAGE ��+`�5TlR~�gQKS~�OFp�KV�0�V_S^]�MPMA2@X_S��$FRCINI�_!U���P�$N)E�P�VTLV�ܠK� �z�%RZ��`b��O2�P�0OV�R10�!�����$ESC_p�uDSBIO�8�`d��.��VIB� �s����e���f��*�SSW.È�VL_���eARM-��Ra���eSC�`�T��Q��MP��rcp�!ru4u5O�ESU�� ��sGwcGw/sGt�s�GtC�Dwɀ'�} �O��IqF��qאSB �F�tG�cgR����7R�v$VOLTt�wN�S�� �� 7Q?T�����PX�ORQF�;���F�?DH_THE@�b�W��a�^�ALPH ^�+�����@ F���N�ɁRM��ӳ��E�p@�3a%2e�1cF�1	M�3aV���Y��9Lr˄INF� �`2bTHR^ <�h�QT԰J�� V=��!t{!o0��1��2 ��{���{�����!�� ���Ӊdd@��ږ��� ���"��1П���"��N��؃CBv�W�IN;HBM�ILT7@=� �d���CP�g�T�����@aaha�da`���@Y�AF��O�઩��� ��ʧ��a`Nô�稧�0R`̩���PL����<#���TMOU���� C������c��CA(�$��?�A̩��I��B��3DI����_�STI�ų۸OX���@����AN���aW$�c0�����$��	���g�_����`RA��`�`fS� ��M�CNUa������V�ERS=��_`I�g�F@��������G�DN4�G.��ǧ�!F�B��ק�M�'�F�_�M>ي � ���Ýt��k֝q�dO2 C��e������DI� ����#� �շ�1���g�Fh ���#�ON�%�a��VAL �CR��_�SIZ��R��1^�REQ_R�|�MBR�|�CHa����ʓ��`|�����*�^�S_E��vh��ggFLG����ge$CV�yM87`�a��FLX@�)B`#bֵe��5AL�`��C_H��T��W����0�b�s � ��NGDMS'�� ��K.c�`_M@X�STW`f� ����AL�` ���a���E���E��IAG�_�to�EJ�T2Ap�� �Q�� �	8p�	Ap�	6�@�_D��!� �
�`��6�Bp=T�� ?�'@!Q.����!L��?O-Y0P.�LD��S�w!�@�FRI�@ �`����A���IV!��NA�UP�`��a��S�LW����`�L-c's'c�C )g��0<���1~���d�a���w(�������"��`�ER�SM� ���F@X$ b�b«tNBAW�q�_TB�m�(PNS_PEA��s�,0���SAV7�(�&WM58��'�CAR��`0�1t4��}2CRQ�� �0�d�3E�P��2STD�ӓ1F�_��7�QOFo��5z%�2RC��6RC˰�86��"Q�bGu 50�gMEA�a_�q���QQآ(�\B~�eDIr�bG�IvbqIgaqG㓣HM���1C�R� ����BF,SDN��Ҏq0��MGqTw1�`�QL ��S�MEf���M�U] !XYZU���A�S�3T>���TRL_@teKX��NU��!U-@�kp+e�pOL*fAR�E��SI�B��E�RWIDT�$�UPP_!P�f1POAW�\E�R���dS7��U* FT�AJN�EMC �~[d(V2_ D_V_h_�_�S`�f3`��P�k�Q�a�U�] ��OV4 )��AN }\C1CRW_I���P��)�h��h�K(�p3�#�X4 P+;�r��?,#v����O��DC��WA2�AOT x$MY� ΃��Xqo�fs�sS�F����D�ҟ����M_SDO��H�LC�����RP��q��C]U?�M17l����`���u>�Z����PNT�V�PL�PV��#��!�p�����@� Pal�1b�BT����vƲ�uNSF�VA�q.S�D	0`Qj���i'5EMA�:�1B�ENY}� ��SUZdۄS�چM�EC)0LD����_����Y�Z�I�I,�I:�#�G.dm�� |��|�,�|�g���H�h����f�EK�PI)d ��K����V�Rβ�CFUNCM�����B�BELW�L��AVI�Bj �t7�� �&)�O��0�TRd�B�A��S��p�r�bS;���A��_DF.�L�� _ 2L ��J��aM��å��`VRl�<���@YLIN���qB�Daߠ�1��H��`MG����EV񑊤THd�4�k�A�1A<�ߣA�EA{�=�1F� �4 RC������`DV���`F����P��	��C�RTP���e 2�Np��cGU���D3NYp��bPK+SA��PK�a�5��ѻGJ�bZDT�2��8��^�DC�%�W�s�c! $���ځ�t%�j#��K@9f������%���0��3C���SW"��EAh��B>�t���B�ACCADJ?�F�p�|1$F��IF4Q�.�JaAF]��?ARGE_Lt���{MOk�$FS�!DS�G@i@z�u���cTPr���`_SJ1 �0�ЛQ{2����4*bY���DIߡ)鄧���J�p�P�AM�Cl/�M�1FU�23s�.�_J5���҃��s�Ct�@CY_ wP LC1IG1h7���J��Mp��2IN�O7��$��CsDEVwICE��Q P2`H�&o��VS���Pfg3�BYl$?�O�PCCs�HNDG7� R� H;�GRP*�E � �b/���Uh����hB��$ CsL�  S0|�g@�b�FB���FEN��&��Cs�X"NqT d2`DO
�PM�9f%^A�K�HOTSW�jDdrV_SELE��Au��~ �BU T82`~�<dNK_x�\�&�[SHA��Z�#$��,�20��'��@7V ���DL��U 
摺��$� �0!;�J$�2�X��3Y{q��T�O:s	&��CsS�LAV�p W � �(�N���Cq_�AR	PUNqX $��CPC_��B �wL'���SH�P�@Y 4�Po��*!�B "?&%?&�R�CF�bZ� 0y�ip#>a�`9f��`�5�aFIL��1�"s��$ID���$� A,��#Wy0�&N�TVt�!V
R�$SKKIZcT�&1<�2�r6J��17 C�06SAF{ �G5_�SV�@�XCLU��Q��2�D_ON�L,�m3Y#=RO=T�HI_VA�Q�PPLY_WARb�3H�P�'�3_Mqv��$:�Y_A.�z�4M��IOC_�1�6CRC1�r�4%3�O됞5LS���$DUMMY47'B A��$} ��y  &3���6|q���cE��XHC����UM��Dర���a���AFsPC	P�#�DTH��pEavP&��NTQ���E,��B�:�s�|"����$TcRY���0�QAs��1_� [ { ��ART_����� �NOC� \�MASTERoԁFYT�!��r!] D��FP_;BA� ��S�!�ђU_^0�\H��S���0��7  ^���cs��If��$!�2]8WSG��� _ � �a�`IGN@�'2a���p��lqh.b%fANN�jGMc��a>�LATCH��`��0rj�g�d�R�.�bDAY�f�U*%` <�q} �#BB�S$��#+C3'H�'A�QEF� I=0 �a @A�ObIT~�"	$TOTA�`*D�A*D	}�EM��NIb��mr�j�nqA�!�t�`���!CAD*�tr+C5r��EFF_AXIJ��c&P�AՃO�p6���N�_R��r!Ed�P�p��Â��Ei���u�PcC�I�MIy��q+� �A8p��qr!e 0�aJ� �yJ��1Z�A ����U@po��CTRLw_CA� f)r�TRAN���IDLE_PWѰ5�F�4IR0V*�V_E��P�e�IAG0Qr!gFw 1$�@| �TKЀ�����0��Pp��R4��ݰAsVE�`����W2�$����9b�u2�Pd���qOH�b��PP2��IRR�	�$BRK��vAB��A��
���R��@� ఐ�*����Pf�x�S@��RQDW�3MS�P��AXe� ���LIFECAL\���L10�N2� ��;�ja0���C��ic{CP�RMOTN��9Y� :aFLA�Cja3OV�aH�HE7a��SUPPO.P���a�]�L= ��ej�_XT_2ʥYӪZӪWӪ�m��>�䣍�_2XZl��Y2.�CO��*�PS�A��N��ja@p��|��P�:RI���o#h `�aACHfSl����ev3m��LA��SUFFIҠ� %���t�rr+C63A�RMSW���i 8��KEYI�MAGMCTM�S��s�"���9a:RO�CVIE<�$qj �BGL�$j`�#�?��P��P�@p#k ��0EN���sm��IN'��B��Mq�B�K�JB�q�q�%ORI_CT�����:a�� ��COF��t�EBU����Pq��	q���q���q����OuF��Hbl ��B�OTh�5�8ң�"0oP_GA�TSCX�����NI_4�j�RО �զ0��I`ICr�O��ճ$�S�ē��M������[�����A(1J`PqiqA��9ӿmL $n�D�o�Io�T�`�$SK�G��$�I�FBK_,�W0DO��RK��@��AW_i�E@p��0��˖@pz�SL����UPCE�B䤯�LE�p_��UF����I�T_�p��Ї�����`��#��>�1_�r�;�2A�1_I7�2Y��qB�n�rT�3T���BUF��՗�~�(��p��PG�o�� xU�y�ղ4 �!@28�p)r}�IR�c��09�o����UP%an�oPm�܄q � ����4�F�5LSP_ ��K�5���s4�1Ë3qE�!dc4�ARR��.�~�T���T�%`�_RD��5���SNeD]�T���VSYP`DZ��2l\���P�m��n-����Po<���� pk���r�R���c+`��~�����Pq ���D�`��s�p$H7OST0!�Pp��	p�4 ��p�EMAIL� ���A�P^�AFAULurtL�}�"�COU� :`;Q�T r!u< �$��%SlЦ�IT�mC��!��DEVI�CE_N�16�SUB��PC�$u��ek!SAVr%4"��M��1F��'�0.5�Py$%ORD=�Q��8X%�A�(OTTp�l�s��@L���*1R�'AX�sp�0X��O3�#�_G2�
PYN_$��%pv�d;FDpp=Dd������F�IF9`�$U�POP7�ED�@EC�`�IwMR�0GH!7q&c�0iqE_aNFOn�x (�PSVv��.t��Iy�rP`wT�y�!��1��#C_RG�IK9bB&b�D]�R4��1}��1D�SP$��2PC`KI cyE�E�1�@U4G��4&�CM�IPV��3p�l�VDTHL�y�GE2�pTJ�WCHS�39C#BSI�[���V�`Z`I�sTy��tNV�@�_G!TL�TF��F�2�5�d9CF�1:aS�C;˕CM��GF�BCMP�S�0ET���z�FU��D�U da��#�WbCD�MI�@� �� �EO�z`}{�s!aI�@�Qe I��!MS���Z�D�Pʔ4�Q) A�|� "�����4�$Z{��NIO#_U<d�{ePàwi�CN��{`l�l�iGROU�W�r���TMN}k u�e u�e p�||�i~cHR�Bp��bw��0CYC{��zsbw~c/⡛zDE�T _D��v�ROpS��qfDAYavq����vTOTz��w�tO4��v�E�4&�AL�0ALa���}�2�!C��!ːBs�i��QRP�%�~~ ,R8�%8�Gz�!LR1} 
�Q]R AUT�2��$������˓$)P�`��C�@��O��5�A1��� H��H *��LX��^` ��VG�P��.���.� �.��.�!�.�.�-�7)�8)�9)�2�+��5�1B�1O�1\�1�i�1v�1��1��1J��2��25�B�2O�U2\�2i�2v�2��U2��2��3��35��3B�O�3\�3i�3�v�3��3��3��4����@�EXT_SEB�Q2��LTЬ��a0w�:e�0FDR�;�T VE	L�#?0	��I⾲�ѷLIFA� +O�VM�ܴA�TR�OV�DT} �M1X���MO�0țIA� ND"�ڲ
Nȋ0?0}�G'1ɱ�`~<1ݱ�� RQ��RI^�MܲGEA-R�IOٵKԲڴ9NF���EFF��P��0qܲZ_MCM�Z`���FEAT�UR�R�y���J!?g ?���? Д?@� �E��(��u4!U�����TP~
q$VARIk��g�4#ETUP2_� � �3#TD�@��2$T�`8ю׈��44"BACK2� QT�4"�4)�:%�PtB�"�IFI`��T��PT�"T�F�LU��}� О�qBGLV�C URS�TYf$�2$P�* �EMP��"$�\�S�?xh�J8��� �#VRTX��0_x$SHO]�L��$ASS�@�C9U�@��BG_��������O���\���i�F�ORCn�p�Kd-��FU�12��2�2j���@"� �|^�NAVYa��\����аS�N�$VISI��s2S�C�$SEFШ�V Oa�$\�а�p�\�$l�I��f��FMR2���F ���Pur���  ����������������Բ_����LIM�IT_
��TC_L�Myƞϰ�DGCL�FY��DY�LD8�|�5��sυ�B0���{�d�'	 T��FS� |� P�S0�3?0$EX_10SP�qj3<5<�G!Qκ�� �^��RSW�[%ONTP
�EBU1G��ٵGR�`a@mUuSBK�aO1��7  PO �P��P{�Mn�O
t`SMo�E�"�@��s`_E � x0� @�TERM%9�%i�ORI�1 Y�%CaSMpOm�B �E&U�M`T(�E&�5�UP�p �g� -?�sb�\��##� �r�G�*� E�LTO�A�p�0<PFI$c�1Ї�P:$�$ߐ$UFR���$���!� �UB OT�7<PT�a��3NS]T�0PAT�q14OPTHJ���PE�P8�3[p�!ARTc �%p� c +2�"RELu:�qSHFT�B�!91�g8_��R�P�SR& ] $l'�0�b����H�c�q�0I�0_U�b} �`PAYLO�@vqDYN_�IЃBp91.�Å�@ERV4� AR�8X�7S�u2��0��_Eߡ��RCH�Å�ASYMFLTR�Å�!WJ�'X�T�E X�c1�IR��QU�DS� Ag5� SF}5P@PC,@Q�6ORS�M��g�GR����	���80� uq��Hm��T�� �?1�֧��POC��!�q$OaP������б,��dbRE�PR�#�qX��a93eB�R75��U�X1��e$PWaR���o�7@R_|S0\4^�t�#UDXӟ3�SVo��PR�" ]�|�$H��!R`�ADDR��H�GP;2ka`aYaTi�Ry��m� Hp�SSC y���eߣ�eO��e\��SE�|�aQRPO}L � � \����bÅ�b�Z�S`UL!LV6tv�_1�V6xj�a��HSCD��O� $H�tP_�p�_�o�MrP?�>��LDT�HTTPu_��Hm� (���OBJ�pYb��$���LE*3�`�q��� � h�+qAB%_O�T��rSEP���,�KR�`�WHIT ����tP��P�r��X�0��P�ןPSS��'��JQUERY_F�LA�!+sWEBS;OC}��HW���!�m��`�@INCPUP^�O���q4�����d���d��\� �IHMI_EDW �T � x��Ht��r�$8�FAV: 4���N��RE��@���@p`E}r�RrQ�Lu��@DFYU3�2$DUMM�Y��H����!IwOLN�Ҟ 8p��R��O�SLR$�INPUT_���$�P��P��#�a�S�LAt �l��������vC��vBT�I�ObpF_AS����$L�Щw�ѹ1�UR �0�!5�r�A�{�@H>���<��MQ��UOP�� ` �Z���2�,�2�3����PP�3�Pz���3���<���P_ME���7� X�IP``Pݢ_NETPe�^�{R������QDSaP��{p���BGP�`a�MaA"� lL"�3TAB�pASPTI���E�� f��0�PSe�BU ID � �Aq���P���a4�L��+0���F�y��Z���Nٸ ڵ�I�RCA_CN� �� ��y��CY�`EA$��w� �x��38�W�RS0�A����ADAY_뀐�NTVA1夰|Ǭ�W5���|�SCA@|�C9L�� ���t��"����X2���N_�PC�����j�=���� �S,ђ��r����fpp� � 3�Q�3���"���c֤rc�LAB+1�� �חUNIH�u�= ICTYs�5�deԂRo �{���q�9�R_U;RL@��$A�`࠰�A^�n g�T�qT�_UW�ABKY_���2DIS\�����iJ��ӡ�ؠ$0∓EyᓀRr�Q�I Aȇ��[�JEqf�FL�%����|�
�wUJR��� ��pF-�7K��'��!����J7��O�B$J�8��7Zo�����7����8���APHMIt�Q�� �D�J7JY�+�*_K�E��  �K�΀LM� � �<��XR�����WATCH_VA��x!@�ѠvFIEL�bVcyi U��խ > b!1V*@Ƶ�CT�и����g �LG��߮� %�LG_SIZ't�� X��FDI  ��� �� �S�� ����. �� ��A{� _0_CM3�,�
��F�A�
���T(���2	/  /��/. ;I.E��/ G9��RS�x�H0  )ZIP�I��0�LN��+R�Zf��DE�E�� ���js�EPL��7DAU�EArp΀hT"	 GHiR����BOO�a��3 C�ѠITW�G$���RE;�^(SC�R�s�DI�S� �`RGI���p�,@����T�"��S�s��W�$���JG=M�'MNCH���FNK��&K7��9�UF'8�0'8FWDv'8HL^9STP':�V'8��'8N '8RS"�9H�@C;�CTt3 �B�Rp�'�9Uiq;4@�'��%��$�.2G9SET?p�y:�%t3��4'�)9EX�TUI5I^ ��^��r�C�#�C0��$	S���	��{%�@z!;NO�FANA�uQ���AI��t���eD�CSm��c-S�c-RO�3XO?WS�]RJXSVX�(IGN ��)01��;�6TDE;a�4LL5!��Ԡi���ñT1$��؜��_�t3A���B����s������+S1%e2%e3%a,�8bB.PԠ� ��{"`T��]%����RqU��?p\&��fST[�R� Y���@�` �$E�fC�k��hp��f�f��Gc�Ԡ� L��*�� ?� ��c�p��h�rpEt���"z#_ �\�ˀ���ļ{ ss�MC��� ��pCLDP|[�C�TRQLI��E�y�tFL,��r����s��D���w�LD8�u�t�uORGK��18�r��ERV��(�Ȼ�(�Ƃ �s��� �耳t�5�t�uv �PT�p��	���>��RCLMC��(�$:���4��1�M���h��b�$DEBUGMAS-�f�W�J�U�$TP��E�����MFRQ~��� � ���HRS_RU���=q.�A<��5FRE�QP!$�  OVER{�)��_f���P01EFI��%�"q/����Q4�U��� \;�h���$U�e`,�?_���P)S$`f�	s�C ���U�����U� �?�( 	��3�IS�C�� d�eaR5Qd�	�TB� ��c \��Ai�AXC��P�l���EXCESH���Q?�M:��Ѽ��aP�C�_�?�SCf`� � H)�`�_�Z�Z�O�񫃯��3�K��Ծߒ�� �B_^��FLICtBh �QUIRE�3MObO�O_�ǖ-�ML?pM�տ mpV!�����=����`MND�x�����!���۳�D��INAUT�!�RSM�����P�N�b��3����ȲPwSTL��� 4��7LOChfRI��he;EX]�ANG	R	�nM�ODA8��L�1�ҧ�~�MF��5 ���i>r�@Hu������SUPDu����FX^�IGGZ! � �_�>s�!� >s�6>t�𹒳bٵ`  ص`/��OC��W��CTI��`�� MN�n�� t��MD��I!)��3P�ԯ���qHq����DIA���a�W�!��a�A��uD#)2�ODO������4 $KHW�NB��N�TIN�aN�#pdI�ǖ��
���`Lk SKªd���Տ�1�_O�q��!sr9 }pT�z�&�Fl��WAI�`O�t�K�EA�����>���V��aL1  � �2T��MpL$ae�|j ��CALL_ጜ�ϑORT�v ���[ ĠCU V��@�y²��� ��T`���^���R_NA �ЈEu��/��U�� OC
TR`�p`�WMp�IA�#����k"4A&PRbS� M�P������ $ F���3�G ǖ�r�!_ꀽ�� ��p0pc���ɒ�����P��� P�KE8�2��$-$B��� ND2��r�2�_TXGtXTRA3S
<��M���ې�P��Yhf���s� SBp�eSWC�SN��M����PU�LS�SNSr�xJ����JOIN� ��p��тr� ?r��p`т��?r��TA&��'P�'�'E�SF�b�RJ~�#ePL$� ư��e�¢D�IR�OB����LO�Aݢ�¢�$� ��&F��e��&�#��M�RR2C��h �6�!_PA���d�E�Ib���G!Q�'2�8<� opRsIN�@ 4<$R0�SW0��M3<�ABC��D_J� V�	����_J3x6
r21#SP��O@	�Pr4�=�3�=j�p	��5JP<��5I��O�QI22��CSKP�zD��$�DJ�A(�QL8EpE8E.Gf�_AZ����1jAEL�Q�2��O�CMPtË�葱R1T ��C�%1�G �%V�`1ͷHY�LZ�D?SMGRST��(�;JGepSCL��a�OSPH_bP(�	U���	�E�RTERpY03�(PA_L�`�Y����P�c(�HTDI܀A�B23U	BDF��jPLWoXVEL��qINSrB�ApB ��T32_��T�W�Wp�UY4Ѓ�0ECH4r<�TSA_Y1�P�GdpT>P��`OFϱ��`��Md`�U*`^�MACC�M��W9 �@�T��E�pв�e�`ep �t_ap_/� �me �bPU���d�"ђi`V�4 DH����� 0 $V
0��S �@[��@~�Y�O��Y��N�RX��H ��$BE`G�(Q_�C`E�QC�3u<�D�IWRC_����T葞��$PS���rL �/su�s�VvF!0@Vv�5y�wKs�w3zr��_1b'���y���5q_MGX�DD��qIRY�FW�ⵂ��Ks6r�DE9�P�PAB)�s��SP�EE�r[�j�IM�.Ar���6qbUS�8�["��P��CTR���Y)�py� ��Y�NB� ȇ�0YɁM�p���pO�P�q��INC�n�8��i�8�31j�ENCY!e�@	�rq6rg�opC�O aIzr_����CNT�S>�UNT23_mRrF��LO~Pr��E.Q D����PGd���a�Fe"��Cx`t�7 I���m �qĂ2CPERC�H  HcO��.R  �t��GѰ�1DGѐG �B����W �3Azrl�L���3��7u��������ƖTRK,U�AY�#f���ۡzr�ߣ�o��FA#�dpMOM�%���Aj�j�T7���'���sq�� DU�20�rS_BCKLSH_Czrm��� ��҂u�?�����0ECLALMq��� ȵCHK
@���GLRTYK��_����$d!����_UM��C%��q�A3Á�7LMT�0_Ln��CL���W�EQ�r�d�P� gum�gx�0���w��ĦP�PC�P�H��MO��CME`C`.�CN_)2N��3Sa@�V����U� (Q��zrV���C� #�SHգ)2�G�$Cc�X��%{q�)�@�PAL"��_P!��_M@�Ub�) 
A����J0	b��\!xPOG׍TORQU���5ޓ���G������G�i�_W4�ۤ�A'���c��T�c��I��I��I�c�F> z��2���1	�VEC5p0���T��1�p����JRK�XH�;���DB�@M�6��MC�0DL�a��GRV����c���c�h�H_3e�����CcOS���@��LNJ� ������@���@����#
��c�Z����h�MY��a������	�THET0��NK�23�c��c��CBֱCB�cC0AS��!�����c��SqB�c�GTSy!��C�1��G���G8 $DU򰏧]P.2�Ul�UQL�_P�(H��CE!KħINX�`�A���3e����LPH������S�## ��/H#2*O�`V�V���`,V*V#+V�1+V?+VM+V[+Vi)H�&2-��%8�#+H1+H?+HM+H�[+Hi)O�O�OT�9.O*O#+O1+UO?+OM+O[+OO�F��-I2D�S�PBALANCE�_q]C`G�p�S�Pea�B�B PFULC�H�B�G�B�Prj1�'�UTOy_��T1T2�I1r2NԱ�r��T!a@&��@��r,s0�T���O�`Nqx�INSE9G�rϑREV6Vϐ�a�DIFǕ�i1�l|W�b1��@OBrQ����B�2qЋ�߱p�?LCHWAR[����AB��D�$ME�CH�q ��Q�AX�P��f��b�@�� 
bf�*qW�ROB �CRzrJe�����C(q_��T �� x $W�EIGH�G�$���c�I偫�IF����LAGւ��S�ւaPւBIL�eO1D�Ґ�bSTBp�bPaQ���`pu�ja
s`�w`
;�(rׁ���  2�ݔ�fDEKBU�cL�p�b\OMMY9ju`PN�ӜKtG�$D�q'��$5p�� 	_�DO_apAra� <�`v�@�ׁ��B�b�`Nq��x_Դ�׀�bOŰ _�� %)�T^��f�9�TsQ-tmpTI�CK�c�PT1up%�sd��N ��@�s �R��ׁ�R��R$�|p_PROMP�E�? $IRI�Ձp��_����MAIm�h��x�_�`v��P��R|�COD�
sFU݀�fID_�����_PY�e@G_SwUFF�� �c4́��DO�VP��`�GR�c�R�� 9���R��R�r����|tpֆ`H�P_F�I	q9n�ORDf�a y`=r36���o�Ձup$ZDT���	E �au��4 *�QL_NA�q�Ȓ�DEF_IؘȒ>��$��b���d��$��>�IS��JДq���W�$���]�;t4ѭ��bDP�@f���
sDF�Og@>�rLOCKE�����*�<�Y����UM ��Ȓ��������e� ������.���f Y�Y���P���Ȓ�@��`�����pP�P G��pS��mpW٨ص�ϣdaTEñ�t��( �aLOM�B_��0�bVI]S ITY�bA�}O�cA_FRI�C�5åPSIS�7��1R��^��^�3#s�bWB:�WF�x�<�L�_���EAS�c��4�P�П�~�_�4\�5\��6�cORMULA�_I����THR.�b��G���w`� �3|8CuCOEFF�_O�qMP`��q!Gd�ѢcS�`\rCA�@�ass$�ác�`�aG�R� � � �$Ϡ$R�rX�pTM§��ϥ�rף�ܦs�ERpPT����h�؛  �BLL���S�_SV��F�#����h��U 5�h�� ���SETUS�MEAn�׀���`�ao�s`�� � ��;` :pг� b�᧡��"͒���á����A��$���D���n�П����P��RE�C���� �pSKy_h@��� P�a?1_USERQ��L�PQL�QVEL@��L�Pt�h��QI����@�MT�qCFG>B��  ��P=O�RNOREq`�p,���SIraߨ�v��RUX����YQͲD�E0 $KE�Y_(s*P$J3OGT`SV7U0a����SW�R=�h����T��GI�@�e`OPWOR� ��,ipSYSsBU� ��SOPu�8���T�
UPPϠ��PAO����R��OP�U�Qؚ�Q��$� IM�AG��*P� ��IM�IN����?RGOVRD� �P��P� �G`b��h��I�RL͠BT�>��PMC_E����9qN�0MxDq=r1�Br��(SL�@C��� � $OVSAL!����,���2�REPq�_(�?�)�@?����=r#C8`�ʐ"#!�)_ZE�R�����$G��� ���B��O @ ?#eORI��"`
}&���)آ!�!��PL����  $FRE�E��E\����PC���t� h� �d���w��PW�R_WS���EN5	1REM8%5	1HWH��3?41сQ9E'!C�� H�a�P��`ATU1SqC_-TDXu6B�Ђ6�k1��}�CqW3��C�� D�q� ���0T�`t�d�"�RXE|0 ���2�2�4r#�y �`�{0UP��o�M�PXb��6�;t3��2� �G���8�SU�Bj1e;�j1�#JMPWAIT@��E�LO>F�qS&RC�VFx�	��R�AREҶ@FWQ�qC& RL��R	��GIGNR_{PL�#DBTB�`PQ��QBW���D��U�p�EIG�H�I��STNLN�F$RR-T[NO��NH�%�PEED@�HA�DOW�`�S��ERVE�vT�8TA�wSPDB�� L�```㑢P��TUN�`�EK�P'AR�0.#LY��@1cbPH_P�KT�$��RETRIE�#����Uk�;FI�"� �y`�P�*d 2��DB�GLV�CLOGS�IZ��KT�AUd>�gdDaS)P_Tc"
��M�C!�&�`vm�R�c���BHEC9KP��L�P��Q�� 0{ h`qAL\� ��NPA��T�R�'t��PIP�#�P��"ARZb���0d�+��\0O��B�ATT �p@+�Zf�`�r��Es�SUXd :"8�� ��Ρ�� $��9IT3CH}B��WO�!��#�qLLB�Q�� $BA)�9D����BAM� U�h��v�!�pJ5 ���r6��q_KN�OW�c�,U��A�D�x�ЭPDO�<�PAYLOA��`�Z��_�1c�xc�Z3L�;�1� L_� !{����q��=��F��C�������I�I��R���~�d�0��B���_J%�!�_J��g��0TAND��?�������!��PL�pAL_� �p�PA��BTk�C��D_�E����J3T�h�� T� PDCKdP�4>��_ALPHx����BEu�2�x�������Qb � �\b�Y�D_1`�2��D��AR54>�(�L�|7��0RTIA4f�u5f�6��MOM��@r����������B�@�ADr��������PUB�R�����@��QAC�h�%��P��"�i�aP���R�q?���� e$PI !=Q�X�e�[�!�*[�Ig�Iu�I��#�@���8A��CA0O��pV# %ZSHIG�s ZS�E�T���T�E�@�@���3���A��A�ESAMP�0�aj���p�8�E�pE� O�� ��M��8@�ƟP)���7�MRO�1m�K0d����KIN��d� S��!��ĚB�G�ԼG�g�GAMM��SX~10rX"ET�"F[ ��D���
$k�I�BRA;RI~AH�I��_�0����E�ސ��A�����LW ��$���H�����t1Pj�C�ECHK64� ����I_R�<p��>��c��ű璣��Ԧ��h� �$�� 1��I>� RCH_DV���aS+�LE��X�!�=����>PMSWsFL�D�SCR-HG100�c`��3nb �����r��ɦ��P���PI3AJ�MET�HO:#���E��AX��#�0X]P��;RESRI��o�3��R�P5�	�$0F��p���IP��B]	L�p�rOOP������APPK�[F�b�`�����RT-g�OS��Pe���2L$�c 1�Z$� ���RA�`MG��!2�SV>���Pp`CURx�LGcRO`P�1c`SA�qcONnbjCNO$0C�! B�j���k� }�������2���(7�DO�QA�ҙa�� ������q�q3�h'�d%"#�� VP�$K$C� S(p� ��!�'p'p � ��S�Ip�&� �Y5�ܐVM_W�RK 2 �%� 0 � �5�!�/8\�/)= )<	L0==`?'p� �N?�?r6�5<<�=�?K1�?�?�OD� BS�;� �1�)� <�?UOgOyO�O�O �O�O�O�O�O	__-_ ?_Q_c_u_�_�_�_�_ �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o �o%7I[m ������� �!�3�E�W�i� Bh�Nc�LMT� l�d9Cl��~�IN������}�PRE_EXEr��ր��_UP갰ʁ1J�!� DV� S�T �'�%?*�J0�Q�HIOOCNV�ȕ��Pl�USʅ5Gi�_�q� 1�+P $��0�v1ϝ�<̟� ?�Z������%�7� I�[�m��������ǯ ٯ����!�3�E�W� i�{�������ÿտ� ����/�A�S�e�w� �ϛϭϿ�������� �+�=�O�a�s߅ߗ� �߻���������'� 9�K�]�o����� ���������#�5�G� Y�k�}����������� ����1CUg y������� 	-?Qcu� ������// )/;/M/_/q/�/�/�/ �/�/�/�/??%?7? I?[?m??�?�?�?�? �?�?�?O!O3OEOWO iO{O�O�O�O�O�M~��LARMRECOV 텰�����LMDG ��Z�-R_IF �����d  YS�T-292 Ma�intenanc�e data d�one se w�ait... R�oot Hub 8Z��_�[pP�_�_�_�o"o0j, 
 �0oYo��8ROS�2 vjLINE �0vaAUTO A�BORTEDvhJ�OIN���o�o�e$�ra  �`�o�m��e�o�\CIO-0�20 LBL[1�] exists� in line� 1:  0 t ew��o�;e	Q�WAYSON_D�O����NGTO�L  � 	 A   ��~��PPINFO 7[ VJ�\�n�����  Cb���� R��ُÏ�����3���W�A�g����@�� ���˟ݟ���%� 7�I�[�m������)��LICATION� ?�u��D`LR �HandHpgTo�olvc 
V9.40P/55�~��
8834�b~�240347��2�������7GDF5�vcN�Q���FRL�� �ub��*�_AC�TIVE�t£�s\���`MODɰ;e��yP_CHGAP�ON����q�OU�PLp1	_Y� �<�@�R�d϶�CU�REQ 1
_[ U �zn�n�	�� ��Ơ��S�ϳ�����������g�1�R;n¤ԥ\��H�u?�r�HTOTHKY��R��\R�d����F� �� $�6�H�Z�l�~��� ���������� �2� D�V�h�z�������
 ������.@R dv����� �*<N`r ���/���/ /&/8/J/\/n/�/�/ �/�/�/�/�/
??"? 4?F?X?j?|?�?�?�? �?�?�?OOO0OBO TOfOxO�O�O�O�O�O �O___,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o0�o�o�o��TO�p˿���DO_CLE�ANϽ�CsNM ; �{ nϑ����t�DSP�DRYRJ��HI�m}@~E�W�i�{� ������ÏՏ�������MAX��*t�a�a�;�X*t:�7�:�>��PLUGG*�+w\7�۵PRC�pBkpEo{4�&���O�����SEGF�K ����k}E�W�i�p{���ş��LAP"� 5�������)�;� M�_�q�����������TOTAL]�3ƟѾ��USENU"��/� xϽb��RGDISPMMC�e��C	�M�@@��/�O �B��+�_�STRING 1���
�M���S��
��_I�TEM1��  n �������������"� 4�F�X�j�|ߎߠ߲�����������I�/O SIGNA�L��Tryout Mode���InpL�Sim�ulated���Out^�OV�ERR� = 1�00��In c�yclR��Prog Aborh����H�Statu�s��	Heart�beat��MH� Faul����Aler�����1��C�U�g�y������� &s��&q�ϲ�  $6HZl~� ������ 82D��WOR��� |��V����� �/"/4/F/X/j/|/��/�/�/�/�/�/�.PO���� 0�	?C? U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcOpuO�O�O2DEV#> �@7?�O�O�O_!_3_ E_W_i_{_�_�_�_�_��_�_�_oo/oAoPALT��ha�Bo �o�o�o�o�o�o�o  2DVhz��p���VoGRI@� ����o�4�F�X�j� |�������ď֏��� ��0�B�T�f�x���R����$���؟� ��� �2�D�V�h�z� ������¯ԯ���
�<���PREGlnU� ȟ.�|�������Ŀֿ �����0�B�T�f��xϊϜϮ���"��$�ARG_|D ?�	������  	�$"�	[�]���"�8���SBN_CONFIG����V�U�o�P�C�II_SAVE � "�x�k���TC�ELLSETUP� �%  O�ME_IO"�"�%?MOV_H���ߎ��REP��!���U�TOBACK����r�FRwA:\B� ,�,B�x�'`��B�u�� �����24/03/�05 00:23�:28B���26 �05:36:02<����52:1��9�B��hꈄA�h�z�`��������B��!`��_D�_\D�02\~W�SLOG.DW�� 2D��`�CRXL.Dkl�������V�  $6HZ�~������ �  ���ATBCKCT�L.TMP CF�G_RPT��PE�AK��_OUTPUT.V�G/Y/k/���X�m�u�>�INIk`��h�|�A�?MESSAG�Ж!�x�С+ODE_D �Ћ�hՉ$�"O�@�/�>�PAUS40 !��� , 	��9��8?F7,		0?j?T?�?x?�? �?�?�?�?�?OOBO�,ONOxM40TSK�  =u�/�A�UgPDT� �'d�@��&XWZD_ENqB�$d��FSTA�%���E��XISV�UONT 2�Fu�w��� 	 �/� rW. ������� �� �ΦB�PP�������u����k_�_�^PQOK  ��kWֿb �i� �#u �ѓ_�_�_�_*on-VMET��2>Y��w�POQA8�y�@��PA 3��?hԱ@?��A&cm>���=v�_>�7��<��+>
P��<��3mSC�RD  1��W� ���u� o�o�o#5Gn� B�9��o����� �S���A�S�e�`w���������$D�GR7P�@�/҃��N5A���	D�φ�_ED� 1�i� 
 �%- EDT-����P�t���˘�:�E�C�B��9�7���<��wp�ܕ2���ß@��D����y���ҟh���ޓ3 ��!���E�W�گE�����4�¯ޓ4}�U�ʿy�2X����X�j� ���ޓ5I����W��r���$�6���Z�ޓ6 ߅�bߩ�W�>ߩ���ߘ�&�ޓ7��Q�.� u�W�
�u����d���Bޓ8�ﹿ��ݿ�X����A����0���ޓ9y�������X���`T�f�����ޑCR� ��R�l�0��TҀ�NO_D�ELޏ��GE_U�NUSE܏�IG�ALLOW 1��}P(*S�YSTEM*z��	$SERV_G�R�z��0REGƚ$�z��NU�M���PMU|=z�LAYI`�z�PMPA�L� %CYC10�1. .W#UL�SU/�3"1��Lm/�$BOXOR=I�CUR_� ��PMCNV&�� 10G.� T4�DLI�@�/�	*�PROGRA�?PG_MI.I?F[0AL)5h?R5[0�B�?�$FLU?I_RESU7'�?���?�4MR�O�
SET��DAT�A-O�$DPMO_SCH���  R�O�O�O�O�O�O�O __+_=_O_a_s_�_ �_�_�_�_�_�_oo�'o9oKo�	ҀLAL_OUT �����WD_ABO�R8 aс�`ITR_RTN  z���j�`NONST�O��d �hCC�FS_UTIL ��ʇCC_A�UXAXIS 3"{ h{ohz���čCE_RIgA_I^�e�p�npFCFG �"}-�!��q_�LIM�2)��Xp� 	��B�\�z���
  �.�z��Zz��N��� ����Y���`��,"�������u�J�z�
3����1����<�#�L�r��PA��0GP 1F|s�����͟ߟ񟰖�CaC��C7�J��]�p������ C���+���+����+���̪��+����+���+���;�� CkT#�+��+��+��+���+��+��+�J���+��+��� D�� D����ڛ��� �޶?��5rHAINFAI�LDO�f)w��EONFI@�o���G_P� 1F{ )Fu(�:�L�^��p���������KPA�US�!1Fu�s G"���Fuܿ� � *�P�6�tφ�lϪϐ� ����������:߰���cA=�u6qM�`N�FO 1���p �1�;����?�?���>Y�L=U��U��Q�C3ҍ�����@��A��;g�`��@����N� ����CD2zD�4��Ca����P��q��4��pO�q ��x~#�LLECT_�ra!���6qM�EN)0p�ei��#�NDER��#�-w1�234567890��Y���r����ЅzByo  )�*�� ��o��H�Z���~� ������������C  2�Vhz�� ����
c.@@R�v���$Z�� g��IO #&�阅N��f-/�?/Q/c/�TR��2'�(����q.��(
-�*�n�_M[OR'A3)F}��� $51�$9<?*?`?N?�?Pr;�"��1*F},�I?������3��K�4���6qP��,Z�� ��-O?OQOɏuO�O�f`�%N�@�܍ON�� �sja�  !}1I�PDB��.�l�cpmidbg�O)_!�;S�:��Up_n_9V/  ��_�_}]܏_[_�_}]/�B�_g�_Doo�^f3o��o,ݑo�ud1�:�o�o{��ADEFg -$�#)�a�c�Qbuf.txAt�o3\�o�0�/�=��>��|2"!6RyMC220�K��d�u�s321�}��t�uN�Cz?���2��BGGA��{�A:L�@$��A"��B����ۮ�_CX�V�B�JA����B�B�C����Q�EŚEM��Dfn6C����D��E�d=�N�>L�͝�Xs6�623�,D>�����!c`2���P�jc`�C
� x��������  D4��C�����  E�%q�F�� E�p��Q�F�P� E��fF�3H ��G�M8��I?��>�3%3~�C���Hn���A�@�B5�\�t2�@At�1�D=x�<#��%�# �O #��-�QzR�SMOFST �+zH�V�P_T1:as4�-A ���MODE 5�=  5���!���A�;�������?����<�M>̼y�TwTEST�b2~��RT�6-���vEC�A݀�H	� Ӂ����r	�C��B��,�C�@���w���:d��# ��Z���Z�r�\�ϡ�T_�`PROG %�:%D��̤ �NUSERi�ѵK�EY_TBL  ��5t����	
��� !"#�$%&'()*+�,-./��:;<=>?@ABC�`�GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~������������������������������������������������������������������������������������������������������������������������������������������[ё�L�CKۼ�Ҵ۰ST�AT!�ͣX|�_A�LM߸���_AU_TO_DO���~v�FDR 38{�2`�AX�q�� EUOSY�ST-325 P�ayload e�rror is �detected� 7920040o1,70��0 ������D$JOGG�ING��1��M�F�AC1��=���B�	i�A?���`�@��Ә"W���Ψ�C@q�C���<{�w�;��� B�P�� B�#��J�@� ��� (Q�}������ C��W���1��CB���B���p�X�R���@��0 Con�tact for�ce excee�ds limit 1,��Y����� ��2G�'�� =�VO�	j�MA?��`���@���c��Z��C��C���$>a���=g+��B�̂��͈�xq��F��� �� ڀ�F���G�����I"�������8��a��s�������G�3�ҧ����@����A�>�`���@��xqf�����CD1�D4��=��77E�B��*��W��b����7� ��� �{�����p2
� �� �o4FX�A�5��{��߂��8���J/���������@W��|���1&�CD22D4�n=&��"�ӣB�� 'B�ȸJ�你�%����oj��Ћ���6��Xz#d��-�?�3G�x?�+*���?�d ���1B�L7�����?��S��l��²��<���fc�B�LC��)D�pA<�V%�2%�JB�; >�AAX�@�.J�m���_����(	�A����+�/?���70�;?M??���O�?�?_�9��5U���1
?Q����v��0�<��y�6�%�C���D�?��ZWSk"B� ݣ���rWO &*�pe+D䘀�_Hxq=��ROdOvO�=��Xze��.�490��4���O�2/co��f�3������=*���(?����ϐA�f�C@���C�<�Cۿc�B�C�b����B������[2:�/�㘀͘�\E��o��̘��'�_*���Xzh�9�O�O_?�CoU`旰VA-� �NK�2߀�A�����ej?���§� ����Af� �]D9�nC���B���d�v��C-���Ђ�M}� [�`����!@���O�"4&5�X{][m�O����O�&��8;S�2��w@j�����3?ܤ�^�K����6���D��C����<�EEw��⵻�B9F_�o���/���a�`/��R����$�/��o�(����e	��p��͏�ߏP�����m <�\7G�5��(���:�@�¡�n�%���c�)��C����C�c�Ct�v�סB��B{�UB>�:h��+����ţ��ᒔ��П���&5�t
��|�-�?���c�u��濙��3G����"���{�@�*¡Z����nc�Y�C��C���Cx|:7�B�P�YB�%'��5-8���@��g��@��3�y�W������{�����1���Ϳ�>߃� <��B��e�@-����yd@S^ ������c�Q�Q�D	YqC�zCw���1ߟ�B������� @��@�� c���ߔ��߸�Rr�tE����_o�b/c�,�����=�<���X=��:�P� �v�O��?���<�ӈ��8�C�G�C濙B=���<\��B�ߊ�b�_�O����$��݃�@��Kx�����CR�� X{^  ���ϟ������9��>h�䊿�~��|*@P�������σ�?�C��I�C朔=Qs[W���Ҽ��o@,��W� ;�`L�T�V�Α��L�P^�p�"9����;�M�_�q�����f	y�{��b��!�W u�7 ������˃�>�C�J/�C�l<����aX�B����bn\��� 1	G����CA�QK���������1CU�/	}�x��� �� v�������?6O �%:#9QY�bB��.@���q*��ŀG�Γ//0/b��5��[/m//�/�/�/�&O	��((� �ys��U�̓�=��O ���R=3�� wB
�B��ݱ��P��K?��@��-N��o��t?(�?�?�����������P_OO�_	����'l��@G������<�C��H1��:>^����Q=t B�~]2�b8YԫO�bAQ����ً�@�A�o��O�O�O�9���%_-_?_�oc_uPJOGGINGMo��o>�G��g���0�� oY@WQ!�����ȃ���'C�/bC濠J=}q7q<H�B�uᇒS."�2=�@��@�	�G�3<�ˑ�O5o�oYo����+{o�o�o`��o�oF��?�S�����3��W n�7 ����u�bC���3p߁=c�5����B���g����O��@��@��kh���G>������.���p�#��5���Y��g�:��� p�wд������
������TC��>�����<�Q����~�Tx[��p���a�"����� �4���4;�M�_�Я������Y�)�ǔ. /k�� �6 <������>~���C���f���>�7��W�m��B���`4�=��f3<�*_��p��p��_�E�PW�ȿ{�����;�������0����f�Y�D�+ǔk��'r� ~�@E����\?��C��C����C曆=@��ڷ���B����Gr�H
o�����N��{q����r�ٿ
X��@�?�?�3�4,70�28>�G�Y����]�P�Ů��#�� {@HUbېR?�����ß��=&�;Ү=�.bB�Lk��%򕰕 W� Ikfxw�� <G��&�8�p�
���\������p��u_&��X?�C'oq��� yH��}ې��=C� O �s@>?-��&w�>�l�B�}gb� A�gw�+ L� F,`�'�S��nqtf7t���

Y� ]������P����9���^���7�� `��@V�ې�_��7@uC�K�C椲<��n��;���B�h�N���U�����9�[9�D�v<�B�f?�(I��� a-�?�cu�9�Ȼ��i��� �8�@IVې�_��7;AC�G�C�U?
6�7!�>�yB� KnGr�߶7 >Hq����G6D3�,`�@,`�/AS j{��?���F?�Y��ף!B�1h��Z���0=��?��� ��9��A�S�C�նC�;��=����1<��nB�G���:OM/���,`n�R��
,`��,~�/�/�/
� m�/�/�/pO�#?5?�OY��cǒ �hv���M�+X?��~��d��J�I�cC���Cؿ��=1�E�A;�X�B��C����rw�? !9�T,`��T�9kaێ�?(OOji o;OMO�_O�_�O�Oo�@��D:�	4��L�>?��7�@ߋ����G2�C��=C��D�=�a8Wa<�ߞB�C�G"���:�?�����9�S n�<禁b�K_]_(o_�/9� Λ_�_��_0�_�_f�A[�g2���A��������y}�#¢nYA�"���B��D;��C��=��B��q<��PBw�A���6��oo�惱��o��o�|�oX�,y�o���C�Ə��m"��p�A������O�y`�¢m�A�#�~�w*D;`�pߌ<�������B���;�	�-������9�_q1��2<�����q�a�"!����%�7�I� W��[�m��🣏U�&���4g2�
��A�f�����E�Yl8��PB'�@�v���DK,OC����=�Q�w�<Կ��B��8��� "/���g�����3���#u�2����!W����͟ߟP���솿ɩG��A��e����M�Y�a.[�2_�b�k�m�DK+�C����>��,ױ=���B���2?Kb���������9�5�#o"�ʯܯ�
��"W���-�?����c�u���)�e�����VA����&���*�G¡�߲BT�Y�C���*DJ��Cֿ
�>� $7�=ׄuB��
��������0� ��S��6<�FU��2�(D�V�(K#W��{ύ���������F�)�i���8A��t���*��*��г��a#ػDJ�C�C�	�=Ď����<���B���%�q=y6
���
�0ܵ�	s����*� �߮��߳�W���������p�#�5����t��g2�QPA�7��3A�-L��м�Z#ֶ��D?ΞC�M��>�����=���{B��~! A�������Q�4����0��w��(����%W��;�M��_��������0����A��2��B�-DDЖ��T����D?���C�T�=	��W{��W{[�W �t2O��vd�0^��:Qn�PTfx�)&W�ț���0/��f/������R8AÐz���.�,�+�¡�Ўa&ӵ�#�D<НCĿ��=)��"�� B��gb=[ �����Z�0%��0��9�0����5�����W�u'W���/&1>/�?M/_/��? �䧲�0��A����9_w�-q� D?��IDD��C�>�YA�=Y5�B���nG҅�.�/�����9`�Q�$W���[D�8?$?6?(�(X�]D[?m?/�Op�?��&_و������CA~}��,��4�����ӿ(�BH�ѣv��LD��C�Q�>Oa�wQ=���B�d�Gҷm�KwO ��) �t��8o�����|O�O��q)�@F�O�O?`Po__�o9Y��GT�A~y]�,�UTWPh[PS_P�cW��D�C�]�>7��a=�zMC"���1/O��+ �D����kƸ�fA�c���_�_�_j��*X�m/o-o�O��co�?�������GR���Au����Ȼ�i��QM�A��I���A�CD���CSLz<Ҩ�17�0��B�ݗ��w7 ���W+ ���3J�+ �gO9���_��+X蒤{������F���0!$���C!Aw�x��i���=Z��A�BA������C�E�CSR�<��엑���{�� @�K*��� ±X��-�$��n�ZB�_��
�|����,X�T{ۏ��?op�#�5����x���rg�1��=�����	i|A?���`�@�������ΈC@�q�C��<t� ��X�Cj�^X�>
���o�?Q�+ ������k�|�OD�-X�qw;��M���п�����D���+�ǣ�=ꫩCӠvנ�۠�ߠ���C@p���!s���*{�T�W� u�"ѮW`��C�U��y����.�����E��5� Payload� error i�s detect�ed 79200�401,70&�8�޿���j��J&Ľ_�=�PӠz7Ϫ颺�.�����5��rA�2M����8G�'��ϵ�q�T��� 
�/�������8/�A�S����}N���=��Ӡ�{נě�δ�Y��ދ�B�M1�����+ ���<��@����9�C8A0��������������&��fǤ�=�ǥ�Ӡ���風�������F�A�u@nq[�v��S���@n�����$��8A1��Ż�����P����CFǤ�=�"@	i�נ�۠�?̙���N5����B���R�!D�[��� ��$�!4����8C�� �$CR_FD�R_CFG 9�?Q?Q��
�UD1:7W�j�$�F&�%s"HIS�T 3:�%#� �   ^xd_Prr� �Q�P_��_*qJ��_F$_nq��_��`_'�$/�_7�M/I?s"INDT_�ENB�S"��.�s"T1_DO0%>Pt5r#T2�?�7�VAR 2;�'.�P t�RE/d��?�|�?d�Z[%��s �STOPi?{2TR�L_DELETE��6 [J_SCR?EEN �%t2kcsc �!�UL@MMENU �1<�I  <xl%xo�O\��O_ (_�b_*_c_:_L_�_ p_�_�_�_�_�_o�_  oMo$o6o�oZolo�o �o�o�o�o�o7  FVh��� ����3�
��i� @�R���v�����現� Џ���S�*�<�b� ��r���џ�����ޟ ��O�&�8���\�n� ������ʯ�گ�9� �"�o�F�X�~���������)�CRE~ =��)�2X�co  ����� A�A7A6JS41�25<@�C_MAN�UALPO{2ZCD�|!>�9�2e� ��"Fn"d���^d�?|(���drǿGRP 2?�9N� B�����?g��� Ҟ��$DBCOb0RIsEs6��G_ERRLOG' @�K!��g��yߋ� �NUM�LIM#1dt5
��PXWORK 1A�KV�������!�3�N=DBTB_�fA BC��#���q���!DB_AW�AY�30  GC;P t2=�׽ҋ�G_AL��d��_ҁYO@sEt0v6��6� �1C�� , 
���� �"�C�M�_�Ma0�!��@�[�OoNTIMpG�t43�}���
����MOTNEND�����RECORD ;2I�K �K�L�G�O�L��� ?Qcu}� �7����F �j�����_ �W/{0/B/T/f/ ��/��//�/�/�/ ?w/,?�/P?�/t?�? �?�??�?=?�?a?O (O:OLO�?pO�?iOO �O�O�O�O]O_�O_H_�NDEXI_�_�_�_�_�_�_�_�NP_C�_$o6o�_ZoEoSo�o�N8}�o�o�oNo ro'�oK]o� �o��8����#��V�TOLER3EN`k�B�����L���CSS_�CCSCB 2J��z��4�L���Ώ ���U��(�:��^�@p���Q�����L���� ����!�3�E�W�i� {�������ïկ��� ��/�A�S�e�w��� ������ѿ����� +�=�O�a�sυϗϩ����� ڟ���L�Y��p�LL{�K����r�P� CL�C���d�L�|�W A�a�pa���������� � 	 3A�����B���?�  ��B�������z��aL�B� L��g��m��ӏ��L������������L���(����@��<:�5�e;��,ȧa���L�Ț ;���x����<����8����\�Ѹ9���>~��:>�+SW��ȝ@��m���>�<,8��?�� Z�����Ȝ��Ad����d�A !Dh�DzuЯ�������W'B(x�_��������K�P�ؐ`0�;C�(  � @��
B�nU�i�oț k�DDȓ>m���C��a����[�YR� ���XZ�ȗ��%/�/I/n/�/�/ȗ�SCHa�t��u�BB�?� D� ?[��/�/ 9/?u��!L�??���2[4J9�Dt4�w29����?!�F1 �3�݈3�7�9�?�? O��?�?OO&OoO�� ��~I0OBO�Oȕ�O �O`��I�/!_3_E_W_ /{_�_l_�_�_�_�_ �_0��dЧ�0hw�\ �om<B��HB�@�X�?�4��r���o55�����>2��;���=ݽw�a� o�o�o�o �R���@Rț�@�@Du�@mx0��@Ed�@��o�B�S�  t�@b�d�!���d�Y�	�d���@��d[� ��@��GY��q�a�1��@j*�d��@��d�Y�ua�d�i�  ��@U��@i�@��@��Y�"�a6�@fa�qY�@|�d��Y��Ъ�b��@��@��d\�C��q2�  ��dF��@%t~�7r�c�Dg�Y�G�b�cF���d��@��@���Y�fT���!��@��d��@�/�d�ۏY�<���*C���d��Y�Q4���F1��d����P��Q��?��������������������C�O¿d�����t�$z��C��h�QA�� A��H A� A��� A�8 A��� A�ɐ؈ �A�� A�  A�0ΐ6��_����H�F72�30-0003-01�*'�9�K�]�o� ��������ɯۯ�����#�5�G��R�0x131EEE70�-{�������ÿ տ�����/�A�S� e�wωϛ��VR������&�  T�S120-602�-1c�/2B3Afb�27�d�C2�g159�/�06M��C�087-901�.�17�93]�o�035}�/�3���� 2���V߈�zߌ�>��v���O������ G����������)�;��M���������u�
��P�
�����6� $Y�y�]
������&8J�ne	o  3�3Մ�#~]pCf�C*� �� Tf�؞)P��C/� ��Q {�P�f��X��\�h����Ä���A�r0>
�@�/%/7/��)nO��vڽ��i�	7U<��ǹ�ߍҼ�"q�' =�U&<�B<��	<��>�&d=ҟ�= Jq<��O�=Yr����=Vy�:*5��;c<���/��O�A*p�/�+O@��?;2Q���Ps0c�B���W�/��O=�=�(A�f#��B����L��f����nA8!��C���A�C���?jO�?�c�	3>�{�ƀA��<`@@�$<`�2�*pBȁ>�3�1C��i`���2�4<��o?�PH�)S�B"p�2,1�1��0�2�B��?5B�
��r��?���b~A�(���0��D`oE�h O�?�OSB���h��?��b�PA(��0�oN�q����S^���X�§lC�9ݪ2�0�A`  ?�0Uo���?��͛4��
m��$DCSS_CLLB2 2OoEo:0<H�u���"y:p�Q8�_�%=0 �n�P�_�?�j�_"o�`��*q� <@�"F�"�� "pA@Ajpce no`�o�o`�@�o�dܖo�d>L9P ��2(3B�?��@An��PD:p@����?�33�aC@~Q�/�RV�@?yC�q��6dw�<a��VV� y�1�AE;� �u��AŴp�u{t� �cu����� a�	���-�?�Q�c� u��������Ϗ�� ���)�;�M�_�q��� ������˟ݟ��� %�7�I�[�m������ ��ǯٯj����!�3� E�W��{�������ÿ տ�����/�A�S� e�wω�߭Ͽ���#��c��TX+1aF#< �߱�aư��� ��o��g��ߝ�K��������=s?�� �_����������C��&LDCKR�EC�Ma�1���)JY���
sF��oIoJ 0���	 ��8\nQ�� �����}���qC �D������� �����/.// R/d/G/�/q/�/ Sew�/*?m/N?`? C?�?g?�?�?�?�?�? �?O�/�/�/\O�/�/ ??�O�?�O�O�O_ "__F_)_j_|___�_ �_5OGO�_�_}Oo�O BoTo7oxo[o�o�o�o �o�o�o�o,>�_ �_F�	o_-o�� #���:��^�p� S���w���ʏM�q ��珹Z�l����� ����Ɵ�����ߟ � 2��V�ُ?�����!� 3�E�����;��.�� R�d�G���k������� ���ǯ��*�<Ͽ�]� 㯄�ǿ�Ϻϝ����� �����%�J�-�n߀� �϶���Kϡ�o�� "�e�F�)�j�|�_�� �����������-� ��T���)��ߜ����� ��������,>! btW����?�� c�u����:}^p S�w���� / �$/�	�l/� %�/	/�/�/�/ ? 2??V?9?z?�?o?�? �?E/W/�?
O�/+O�/ ROdOGO�OkO�O�O�O �O�O�O_�O<_N_�? �?V_�_Oo_=O�_�_ 3_o�_%oJo-ono�o co�o�o�o�o]_�o�_ "�_�o�_j|�o� �������0� B�%�f��oO��1 CU���K�,�>�!� b�t�W���{���Ο�� ��׏��:�L�Ϗm� 󏔯ן��ʯ��� � �$��5�Z�=�~��� �%�ƿؿ[���� � 2�u�V�9�zό�oϰ� �ϥ�����
�ߟ�=� �d��9�Ϭ߾�� ���������<�N�1� r��g��+ߑ�O��� s߅ߗ���J���n��� c������������� ��4�����|��� #�5����0 B%fI��� �Ug//�;/� b/t/W/�/{/�/�/�/ �/?�/(??L?^?� �f?�?)/?M/�? O C?$OO5OZO=O~O�O sO�O�O�O�Om?_�? 2_�?_�?z_�_�O�_ �_�_�_�_
oo�_@o Ro5ovo�O___�oA_ S_e_�o[o<N1 r�g����� ���o�oJ�\��o}� �����ڏ����� �4��E�j�M����� #�5�֟�k�����0� B���f�I�������� ү����ٯ�,���M� �t���I����ο� ���(��L�^�A� �ϔ�wϸ�;���_� � �������Zߝ�~ߐ� sߴߗ�������� � �D���)��`�V�� �������������8�7�I��>l����2k�  ������{������ ��������FXj� g�C(  @�@  A�Ӈ@��{A   ?���?�� � g�@���ffC�!�	� Bp� �  �F?����@�l#��   �B� B�  C�J�� `!�UHf�� �A 5�L�� �������	� � A� ��� ��$DCSS_C�NSTCY 2P����  md����/ /4/B/T/f/|/�/�/ �/�/�/�/�/??,?�>?�DEVICE 2Q�#�5"�&�T?_��?�?�?�? �?OO(OUOLO^O�O �O�O�O�O�O�O	__�-_�F�HNDGDg R�$�Cz���LS 2S� �_�_�_�_�_�_o�o:_�PARAM7 T��bT���Q�2�RBT 2�V� 8 
 <�?} � ���� �E�R�8�lʹa��0�W  �eB\�o�f���MCp�%.w#���o�f>�K0�����q$��n� �逨f���|�b�u���FcRj� ��]�4��F�e�j�|����IC���DjPC�$Z���@���A,���4�u@�X�@��^@w��|�J����B��%��C4�C3:^C4���A����8�-�B{B���A���&�l���C�C3��JC4jC3���d� +�3 D�ff 2�A PЩ��K@�d����� ��ן�����l�C� U���y���������ӯ  ���	�V�-�?�Q�c� u���Կ����
�ϗ� 4�F�1�j�Uώ�yϲ������� ğ��ڿ ��g�>�Pߝ�t߆� �ߪ߼�������Q� (�:�L�^�p����� ������� �M���q� \��������������� ���.�#�DV �z������ �
W.@�dv ����/��A/ /*/I/�/�/�/�/ �/�/�/�/+??O?* X/j/�?R/�?�?�?�? �?O�?�?KO"O4OFO XOjO|O�O�O�O�O�O �O�O__0_}_T_f_ �_�_@?�_�_o�_1o oUo@oRo�of?�_�_ �o�o�o	�o�o (:�^p��� ����;��$�q� H�Z�l�~������jo ��%��I�4�m�X��� |���ǟ�oЏ��� ��E��.�M�R�d�v� ï������Я��� �*�w�N�`������� ����̿޿+Ϧ�O�:� _υ�pϩϔ��ϸ��� ̟ޟ�����"�4߁� X�j߷ߎߠ߲����� ��5���k�B�T�f� x������������ ��g��ϋ�v������������	��-:	��$DCSS_SL�AVE W����[�~D
_4D  [�pAR_MENU X[ "�� ��6��@�R@�SHOW �2Y[ �  /?��������/"/(F/X/j/  ��/��/�/�/�/�/ ?4/1?C?U?|/v?�/ �?�?�?�?�?�??O -O?Of?`O�?�O�O�O �O�O�OO__)_PO J_tOq_�_�_�_�_�_ �O�_oo:_4o^_[o moo�o�o�o�_�o�o �o$oHoEWi{ ���o@��, 2/�A�S�e�w����� ���я����+� =�O�a�s��������� ������'�9�K� ]�o���������ޟد ����#�5�G�Y��� }�����ȯ¿���� ��1�C�j�g�yϋ� ����ֿ������	�� -�T�Q�c�uߜϖ��� ����������>�;� M�_�߀�ߧ���� �����(��7�I�p� j������������������!3eCFG7 Z{�������FRA�:\sL}%04_d.CSV@	 m}@ �A �CH� zd��[�����h�.�@R��JP��n2  �ASRC_OUoT [^h���_C_FS�I ?� �&//// X/S/e/w/�/�/�/�/ �/�/�/?0?+?=?O? x?s?�?�?�?�?�?�? OOO'OPOKO]OoO �O�O�O�O�O�O�O�O (_#_5_G_p_k_}_�_ �_�_�_�_ o�_oo HoCoUogo�o�o�o�o �o�o�o�o -? hcu����� ����@�;�M�_� ��������Џˏݏ� ��%�7�`�[�m�� ������ǟ����� 8�3�E�W���{����� ȯïկ����/� X�S�e�w��������� �����0�+�=�O� x�sυϗ��ϻ����� ���'�P�K�]�o� �ߓߥ߷��������� (�#�5�G�p�k�}�� ������� ����� H�C�U�g��������� �������� -? hcu����� ��@;M_ �������� //%/7/`/[/m// �/�/�/�/�/�/�/? 8?3?E?W?�?{?�?�? �?�?�?�?OOO/O XOSOeOwO�O�O�O�O �O�O�O_0_+_=_O_ x_s_�_�_�_�_�_�_ ooo'oPoKo]ooo �o�o�o�o�o�o�o�o (#5Gpk}� ���� ���� H�C�U�g��������� ؏ӏ��� ��-�?� h�c�u���������ϟ �����@�;�M�_� ��������Я˯ݯ﯀��%�7�`�[�m���$DCS_C_F�SO ?������ P s�m���߿ڿ ���'�"�4�F�o�j� |ώϷϲ��������� ��G�B�T�fߏߊ� �߮����������� ,�>�g�b�t���� ����������?�:� L�^������������� ����$6_Z l~������ �72DVz ������/
/ /./W/R/d/v/�/�/��/�/�/�/�/�C_RPI����
?S? |?w?"?��F?�?�?�?,�?��SL4?@�?O QOzOuO�O�O�O�O�O �O
___)_R_M___ q_�_�_�_�_�_�_�_ o*o%o7oIoromoo �o�o�o�o�o�o !JEWi��� �����"��/� A�j�e�w��������� я������B�=�O� a���������ҟ͟ߟ ��� O�?DO&�o� ���������ۯ��� (�#�5�G�p�k�}��� ����ſ׿ ����� H�C�U�gϐϋϝϯ� �������� ��-�?� h�c�u߇߽߰߫��� ������@�;�M�_� ������������� ��%�7�`�[�m�� ���������������83�<NOCOD�E \�5���;PRE_C�HK ^�;J A� J �<� �O �5���5 	 <�W�� =O)s�_q� ���/�'/9// %/o/�/[/�/�/�/�/ �/��/#?5?�/Y?k? E?w?�?{?�?�?�?�? OO�?+OUO/OAO�O �OwO�O�O�O�O	_�/ ??_Q_�O]_�_a_s_ �_�_�_�_o�_o;o o'oqo�o]o�o�o�o �o�o�o�o%7[ m'_U����� ��!���W�i�C� ����y�ÏՏ����� ���A�S�-�w��� q���џk������ =��)�s���_����� ��ǯ�˯ݯ'�9�� ]�o�I�{�������ۿ ����#����Y�k� EϏϡ�{ϭ��ϱ��� ����C�U�/�aߋ� e�w����߭���	�ÿ ��?�Q�+�u��a�� ���������)�;� �_�q�K�]������� ������%�[ m��}��� �!�EW1c �gy����/ �/A/7Iw/�/#/ �/�/�/�/�/?�/+? =??I?s?M?_?�?�? �?�?�?�?�?'OOO ]OoOIO�O�O_/�O�O �O�O_#_�OG_Y_3_ E_�_�_{_�_�_�_�_ o�_�_CoUo/oyo�o eo�o�o�O�o�o	�o -?KuOa� ������)�� �_�q�K��������� ݏ�o�o�%���1�[� 5�G�����}�ǟٟ�� �����E�W�1�{� ��g���ï������� �/�A���)�w���c� ���������Ͽ�+� =��a�s�Mϗϩσ� ���������'��K� ]�S�Eߓߥ�?����� ���������G�Y�3� }��i�������� ���1�C��O�y�o� �߯���[��������� -?cuO�� �����) 5_9K���� ����/%/�I/[/ 5//�/k/}/�/�/�/ �/?�/3?E??1?{? �?g?�?�?�?�?�?� �?/OAO�?eOwOQO�O �O�O�O�O�O�O_+_ _7_a_;_M_�_�_�_ �_�_�_�_oOOKo ]o�_io�omoo�o�o �o�o�oG!3 }�i����� ��1�C��g�y�3o a����������я� -���c�u�O����� ��ϟ៻�͟�)�� M�_�9�������}�˯ ݯw�����I�#� 5����k���ǿ��ӿ ��׿�3�E��i�{� Uχϱϧ������ϓ� �/�	��e�w�Qߛ� �߇߹��߽����+� �O�a�;�m��q�� �����������K� ]�7�����m������� ������5G!k }Wi����� �1'�gy �������/ -//Q/c/=/o/�/s/ �/�/�/�/??�/#? M?CU�?�?/?�?�? �?�?OO�?7OIO#O UOOYOkO�O�O�O�O �O�O	_3___i_{_����$DCS_�SGN _k5��%)���18-JUL�-24 12:1�0 ]S05-�MAR�Q00:4�1�P�P�R �XzaE�RehXeU�Q�R�Y�P��Q�RB,�Þ����E��_�P�o���5���X��K�_U~�THOW `k5 �Q��UVERSION� �V�`�?V4.5.8�Y�P�EFLOGIC �1aui�  	\Pfp0�ip0�n�b�PROG_ENB  �T�c�P	sULSE  �e�!u�b_ACCL{IM4v�#s�dHsWRSTJN�T4w�a��TEM�O|�Q%q�b�pINIT b�jg:�`��tOPT_SL �?	k6�r
 	�R575�S�p7�4�y6�x7�w50
�1�2�t�hG��g>�tTO  �}#ot���fV�pDEX4w�d�b�P��PAT�H A�jA
\�18072024�\ UME IN�FORMAT�`\�����cHCP_CLNTID ?�f�c �h�UR���bIAG_GRP� 2gk5a���R	 @��  ��ff?a�G����Z��B�  ȟ�\ő�ΐ�ߞ�@c���!�7�@�z�@^��@
�!�Ym�p3m29 89�01234567�E��ws0� ����Rd�h�}��Va��Q�B4�����X  �U�xͣa�_�k6�� �>�k6Ѡc>�������-�ǿQ�c�u��\�ԿϨ���T�޿ �ϜϮ�8϶���n� �ϒ�,�>���b�t��� l�xߺ�Dߪ����� ��8�J�(�Z��
�� f�����������4��q2c�d�!� Ѹ�?��x�@`�������5!���4V�ɕ����A�P��@�����Z��?�����������8�F�=q��=b��=�E1�>�J�>�n��>��H��<�o� D
�sT�\�N���QCp  <w(�U�R 4��i������YA@�R?���@��� i8�F�V|^x��D�>J����bN�����Gy����@���$"�?��0!/@ff�!6 M!�33�X"(��޸�C�� t"I���CH�)C.dBت��΢�/�!�,'6p�/��͐�%�B�P�%d.[ 1B���7�/=?O?B XT��G�	���P�?���>&�?\��?����܁>��M��.J�����CD2LD4�� �P(���Q?�?�?�?�(��?BR9�9C�a~���+�?�K<�&`�?QO �?uO`O�O�O�O�O�C�:=�_����B���ة�;D{��U:�oU�n�CT_CONF_IG h���s>�Teg�ez��STBF_TTS4w
!yhS�`4s�Q{Vh`MAUop�b�MSW_CF<Pi  �lOCV7IEW�Pj�]Ñ��g�!o3oEoWoio {oMRo�o�o�o�o�o �o�o"4FXj| ������� �0�B�T�f�x���� ����ҏ������,� >�P�b�t�����'��� Ο�������:�L�`^�p�����$\PM�R�k�]RSͧШ
� έ����SC�H 2r�[
|�ScheduOle 18k oRQ`
R4��`��*3�ϥ��]�R;��MQ>L�ͯ���ܿ���� ˿$����l�7�I� [ϴ�ϑϣ������� ��D��!�3ߌ�W�i�p{��ߟ߱�	 l�������PST�`	�� R9Dz.����#�5� G�Y�k�}������ ��������1�C�U� g�y������������� ��	-?Qcu ��������);M�NR5= ��������//)/;/M/_/q*	���/ �/�/��I VB�T�? x���K?�߸�:?�?^? p?�?�?�?�?�?#O�?  OOkO6OHOZO�O~O �O�O�O�O�O�OC__  _2_�_V_ �r�� ��`�_�_�_�_
o o.o@oRodovo�o�o �o�o�o�o�o* <N`r���� �����&�8�J� \�n���������ȏڏ ����~/|/���� ԟ���
���/L�^�p��/�"%�21��/? �)?{_��_i_�`� +�=�O���s������ ��Ϳ߿8���'π� K�]�o��ϓϥϷ�� ������X�#߱_#�5� G�Y�k���ߡ߳��� ��������1�C�U� g�y���������� ��	��-�?�Q�c�u� �������������� );M_q�� ���}�/�Yk} �����1�C�/ +/=/���/˯�/�A� �/e�/߱/
?�/�/�/ R??/?A?�?e?w?�? �?�?�?�?*O�?OO rO=OOOaO�O�O�O�O _�Ow���1 �_9_K_]_o_�_�_�_ �_�_�_�_joo#o5o GoYo�o}o�o�o�o�o B�o�o1�U gy������ �	���-�?�Q�c�u� �U��'�9�K�]� o�����	/ß՟�Q/����3��o/�/^��/ �O��_�O��ܯ���� ˯$����l�7�I� [����������ǿٿ �D��!�3ό�W�i� {��ϟ�-_����ÏՏ 珍���/�A�S�e� w߉ߛ߭߿������� ��+�=�O�a�s�� ������������ '�9�K�]�o������� ����������#5 G������� /AS������� �i/G�/k���>/�� ��-/�/Q/c/u/�/�/ �/�/?�/�/?^?)? ;?M?�?q?�?�?�?�? �?�?6OOO%O~OIO ��ew���_�O �O�O�O�Oz_!_3_E_ W_i_�_�_�_�_�_�_ Ro�_oo/oAo�oeo wo�o�o�o*�o�o�o �=Oas� ������n�� o������Ǐُ��� ��?�Q�c���%�4)���ڟ!/sO� �OaO��X�#�5�G��� k�}���诳�ůׯ0� ����x�C�U�g��� �������ӿ���P� ϩO�-�?�Q�c�	� �ϙϫϽ�������� �)�;�M�_�q߃ߕ� �߹���������%� 7�I�[�m����� ���������!�3�E� W�i�{���������u� '�Qcu���� �)�;�#5��� ß��9Ϻ]�'ϩ /���J//'/9/ �/]/o/�/�/�/�/�/ "?�/�/?j?5?G?Y? �?}?�?�?�?�?o��� ��)�O1OCOUO gOyO�O�O�O�O�O�O b_	__-_?_Q_�_u_ �_�_�_�_:o�_�_o o)o�oMo_oqo�o�o �o�o�o�o~% 7I[m�M�� �1�C�U�g�y���@��͏ߏI����5�� gyV���?��O�? {�ԟ����ß���� �d�/�A�S���w��� ������ѯ�<��� +���O�a�s�̿��%O �������� '�9�K�]�oρϓϥ� �����������#�5� G�Y�k�}ߏߡ߳��� ��������1�C�U� g�y���������� ��	��-�?������ ����'9K�� �������a?�  c���6ٿ��%~I [m����/� ��V/!/3/E/�/i/ {/�/�/�/�/�/.?�/ ??v?A?�]�o��� ����O�?�?�?�?�? rOO+O=OOOaO�O�O �O�O�O�OJ_�O__ '_9_�_]_o_�_�_�_ "o�_�_�_�_o�o5o GoYoko}o�o�o�o�o �o�of��g��� �����}7�I�[����6!��� ҏk?��?Y?��P� �-�?���c�u����� ����ϟ(����p� ;�M�_��������� � ˯ݯ�H���?% 7I[������� ǿٿ����!�3�E� W�i�{ύϟϱ����� ������/�A�S�e� w߉ߛ߭߿������� ��+�=�O�a�s�� ����m�I�[�m� ���������!�3�	 -{����|ߏ1� �U������� B1�Ugy ����/��	/ b/-/?/Q/�/u/�/�/ �/�/g��������!� �?)?;?M?_?q?�?�? �?�?�?�?ZOOO%O 7OIO�OmOO�O�O�O 2_�O�O�O_!_�_E_ W_i_{_�_
o�_�_�_ �_�_voo/oAoSoeo �oE���);M _q������A����7��_qN�� �/��?�/s�̏���� ���ߏ��\�'�9� K���o�����쟷�ɟ ۟4����#�|�G�Y� k�į��?�o�o�o�o �o}o����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� �)�;�M�_�q߃ߕ� �߹���������%� 7��o���������� �1�C��������� �Y7���[���.ѯ ��vASe�� �����N +=�as��� ��&/�//n/9/ �U�g�y����/�/ �/�/�/�/j??#?5? G?Y?�?}?�?�?�?�? BO�?�?OO1O�OUO gOyO�O�O_�O�O�O �O	_�_-_?_Q_c_u_ �_�_�_�_�_�_^o�� _��o�o�o�o�o�o�o �ou�/AS����8������c/ � �/Q/�H��%�7��� [�m��؏����Ǐ � ����h�3�E�W��� {�������ß՟�@� ��/oo/oAoSo�_ w���������ѯ��� ��+�=�O�a�s��� ������Ϳ߿��� '�9�K�]�oρϓϥ� �����������#�5� G�Y�k�}ߏߡ߳�eo A�S�e�w���� ��+��%�s�� �t��)���M���� ��������:) �M_q���� ��Z%7I �m���_��� ������z/!/3/E/ W/i/�/�/�/�/�/�/ R?�/??/?A?�?e? w?�?�?�?*O�?�?�? OO�O=OOOaOsO�O _�O�O�O�O�On__ '_9_K_]_�_=����_ o!o3oEoWoio{o��@�o�o�o9��p9� W�i�F���|/� k������� �T��1�C���g�y� ��䏯���ӏ,���	� �t�?�Q�c�����/ �_�_�_�_�_u_�� �)�;�M�_�q����� ����˯ݯ���%� 7�I�[�m�������� ǿٿ����!�3�E� W�i�{ύϟϱ����� ������/��_�o�� ��������)�;�o �o}����oQ�/�� S��&�ɟ���n�9� K�]������������� ����F#5�Y k}����� �f1۟M�_�q� �ߕ������� b/	//-/?/Q/�/u/ �/�/�/�/:?�/�/? ?)?�?M?_?q?�?�? O�?�?�?�?O~O%O 7OIO[OmO�O�O�O�O �O�OV_��W�y_�_�_ �_�_�_�_�_m�'o9ohKo���hv10w ��o�T�oxB �o9(�L^ p�������  �Y�$�6�H���l�~� ��鏴�Ə؏1���� �_ _.�D_���Oz� ������-�ԟ���
� ���@�R�d�v���� ����Я���q��*� <�N�`�ݿ�������� ̿I����&�8ϵ� \�nπϒϤ�!�h_o D�V�h�zߌߞ߰��� o����do��o�o w��oh��P����� ����������,�>� P�b�t����������� ����(:L^ p����b����� ��
����$6HZ l~������ �/ /2/D/V/h/z/ �/�/�/�/�/�/�/
? ?.?@?R?d?v?�?�? �?�?�?�?�?OO*O <ONO`O.����O __ $_6_H_Z_l_��$�_��_*�<��$DRC_CFG sE�?�!L�o �JoKo:ooo^o�o�o��o��PSBL_FAULT t	j��e�dGPMSK � �d�g�PTDI�AG uE�gQ�P����UD1: 6�78901234�5Ar�5q\��P �o����� ���!�3�E�W�i�@{����oY�4s��@�C�m��eTRECP,z
:t,�Sw/�k h�z�������ԟ� ��
��.�@�R�d�v��������ӏЯ�gUM�P_OPTION�`�n�TRb�c�i=�PMES�	��Y_TEMP  È�3B�� �_��A\�I�UNI�T�g_�vYN_B_RK v	�(r~��EDITOR����8���_�ENT� 1w	i�@,&�ROS2  O�Rr����J&PR�OVA��2�&	?TRANSP"�4�&DE�c{�
Χo������������ ���5��Y�@�}ߏ� v߳ߚ���������� 1��*�g�N��r�� �������	���?��&���MGDI_SCTAr��_�� ���NC_INFO �1x���������3����~�f�1y�� ������� �E d��M_q� ������ %7I[m�� �����//") :"/H/Z/l/~/�/�/ �/�/�/�/�/? ?2? D?V?h?z?�?�?�?** ��?�?OO1/;OMO _OqO�O�O�O�O�O�O �O__%_7_I_[_m_ _�_�_�_�?�_�_�_ o)O3oEoWoio{o�o �o�o�o�o�o�o /ASew��� �_����!o�=� O�a�s���������͏ ߏ���'�9�K�]� o���������۟� ����+�5�G�Y�k�}� ������ůׯ���� �1�C�U�g�y����� ��ɟӿ���	�#�-� ?�Q�c�uχϙϫϽ� ��������)�;�M� _�q߃ߕߧ������� ����%�7�I�[�m� ������������ �!�3�E�W�i�{��� ������������� /ASew��� ����+= Oas������ ��'/9/K/]/ o/�/�/�/�/�/�/�/ �/?#?5?G?Y?k?}? �?���?�?�?�?/ O1OCOUOgOyO�O�O �O�O�O�O�O	__-_ ?_Q_c_u_�_O�?�_ �_�_�_Oo)o;oMo _oqo�o�o�o�o�o�o �o%7I[m ��_����o �!�3�E�W�i�{��� ����ÏՏ����� /�A�S�e�w������ ��џ����+�=� O�a�s���������ͯ ߯���'�9�K�]� o���������ɿۿ�� ��#�5�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߓ��� ����������	��-� ?�Q�c�u����� ��������)�;�M� _�q����ߧ������� ��%7I[m ������� !3EWi{�� �������// //A/S/e/w/�/�/�/ �/�/�/�/??+?=? O?a?s?�?�?�?�? ��OO'O9OKO]O oO�O�O�O�O�O�O�O �O_#_5_G_Y_k_�? �?�_�_�_�_�?�_o o1oCoUogoyo�o�o �o�o�o�o�o	- ?Qc�_�_��� ��_���)�;�M� _�q���������ˏݏ ���%�7�I�[�m� �������ǟ���� �!�3�E�W�i�{��� ����ïկ����� /�A�S�e��m����� ��ٟϿ����+�=� O�a�sυϗϩϻ��� ������'�9�K�]� w����ߥ߷�m���� ���#�5�G�Y�k�}� ������������� �1�C�U�o߁ߋ��� ����������	- ?Qcu���� ���);M _y�������� �//%/7/I/[/m/ /�/�/�/�/�/�/�/ ?!?3?E?W?q{?�? �?�?��?�?�?OO /OAOSOeOwO�O�O�O �O�O�O�O__+_=_ O_i?[_�_�_�_�?�? �_�_oo'o9oKo]o oo�o�o�o�o�o�o�o �o#5Ga_s_} ����_���� �1�C�U�g�y����� ����ӏ���	��-� ?��ku�������� ϟ����)�;�M� _�q���������˯ݯ ���%�7�I�c�m� �������ǿٿ��� �!�3�E�W�i�{ύ� �ϱ����������� /�A�[�I�w߉ߛߵ� ����������+�=� O�a�s�������������'�9�S� ��$ENETMO�DE 1z���  cЅc�^Հ���b�O�ATCFG {^���������C���DATAW 1|o����**��1HCUddd��� ����k����Zl~����7I�//,/�P/�����/@�/�/�/?/�/��o/ �/.?@?R?d?�/�?��??�?�?�? Ow?$O���?�?fOxO�O�OO�OZ�RPOS/T_LO��~��^Ձ
��	__-_?_�BR�OR_PR�@%�o�%]�x_G_R_TABLE  o�����_�_�_�WSRSEV_NUM ~�4�y�`�A�_AUTO_EN�B  ��w��D_;NO-a o���}b  *�p`��p`�p`�p`#`+�o`�o�o�oIdFLT9R5oGfHISc2�@m_ALM 1��o� �g%pl]�+�oI[m��r�o_bO`  o��na���zb�TCP_VER !o�y!p_�$EXT�@o_REQ�f�@i�:�SIZC�5�ST�K`�^e�7�T�OL  `�Dz��b�A 5�_BWD�p���fɁ��;DI�� ����Gx��ϊSTEPߏ��b��OP_DO���`�FDR_GR�P 1�o��ad �	�����q�s��V��'�N"����l��?T� �����q� Ɵם������	�B��-���_>���8��s������>�׽E��T,���P���ï��<���>?�z@�;3�@	��>���hܡǪ
 K�Zw`��l�ǯv��ȯ��W�B�{��f�A@  ��@S33��`�@����_�x���q�F@ ϼռq�G�  8�Fg�fC�8RDŞؽ?�  `���6��X����875�t��5���5�`+�ؽ��t���[JW��Ǖ8�0��p���KFEATURE ����ɀ��LR� Handlin?gTool �`��Englis�h Dictio�nary�4D ;St��ard���Analog I�/O6�?�gle �ShiftR�ut�o Softwa�re Updat�ew�matic ?Backup٥��ground E�dit���Cam�eraM�FQ�Co�mmon cal�ib UI����n�����Monito�r �tr �Rel�iabf��DHC�P���Data ?Acquis�8�?iagnos��J�~R�isplay��?Licens6�<��ocument �Viewe�:�u�al Check Safety��~�hanced��4���s��Fr����xt. DIO ��fi���end.��Err�L��8�J�s7�rH�'� ����FCTN Me�nu��v6��TPw Iny�fac���GigE�������p Mask Ekxc��g�HT���Proxy Sv�����igh-Spe��Ski������~+�mmunic��7ons2ur��y��M�Nѳ�conne�ct 2incr��stru�g
� �e����J���KA�REL Cmd.� L��ua���R�un-Ti�Enyv�z�el +��s��S/Wע������N�Book(S�ystem)�M�ACROs,)/�Offsem�LH0+���K�QMR�⢆�M��| *�l��MechStopt� l�LiI�i��ax��JТ�{odg�witch/�{�y.q,+Optm>/L� fi��g_~Lulti-T������PCM fu�n��)a�tiz��(�'oi�Regi�ArM �&ri��F��+6K�Num S�el�'9� Ad�ju= ">O1i�`=t�atu1x?���R�DM Robot>�scoveѴ5�ea� �Freq� AnlyMRe�m�+�n-״5�2S�ervo+� �S�NPX b	n�SN��Cli��7NjҏLibr�WO�� ��i@#Fo&t��sGsag�%�D�p Әd9��p/I���EM�ILIB�O�BP OFirm���NP���Acc����TPT9XG�Delnd�O�A��`�Morqu>g�imula���tVu  Pa�N��t4�:#& ev.�E��ri��L_US?R EVNT�_`nexcept����0n�� e�S�VC"��rH?�Vh�eb�_veiKpkSJ@SC�FU�oSGE�o�eU�I9�Web Pl �6�nA_t ����n�ZDT App�lF�WqEOATX�A���iPB�aPI>� Grid�1��\�}|iR\b.-���v{�}o��RX-1�0iA/L�Al�l Smooth�-��s�S���Pri�tyAvoidM
�s/�t�P?���V01o���!��ycf��00�P��;�CS� g. c�⼈Jo1 � ф׏$҂����M�t|��c�abo�4~��main N�A.8�yp y� isfi����PMC����RL�P�
y��av����p��bc���MI Dev�� �(+AE�y�d�1/ ��ַS��"�1��0iC�rt(�en��4��ni+��!<���'sswo4���ROS Eth
��P��eMw�4�9L�X� b���E<�Up0N0A�E3�t ���Wr0 down�-al�Puero D N��V ��z�
v�v�K4��8�64MB �DRAM4���FR�O��}�X�� Fl�  �0`�� r�2�o�s�n�Ce8�N���shD�P�b�c]+_Ņ�Yp�Vt�tyf�s92 ����ᯧ��2V _���́/s���d��0Xk�O�� 2��a|��por*�EMAILB{~�Q���MK��h�0B.�q��T1�cFChe��Fs莿�Hel�u�޿3T[yp��FC h��t��*`SLFor��(�r�lu �42��LCMGRH_NP'G j�}R�zz/��1reP0)�Net�Fr)г���o m��0�0c���tOPC'-UA��3�T1�� dA���S�p��cr�v�+lu�@ AP�e ����!(7( �3�t��:�Qp�PSyn.�(RSS)�6quires �@'��3�iE�tN���est~�EIMPLE ��f"G��LM#FS��e�Btex�T��!H�plQ3b�_CPP �ExO�?+��`x�Tea  tY���Vɠ��#ru�&(�!S��Q��xۑ��@�fUIF�ƒoni��ustdpn�[�t��r�� ����+/"/4/F/ X/�/|/�/�/�/�/�/ �/�/'??0?B?T?�? x?�?�?�?�?�?�?�? #OO,O>OPO}OtO�O �O�O�O�O�O�O__ (_:_L_y_p_�_�_�_ �_�_�_�_oo$o6o Houolo~o�o�o�o�o �o�o 2Dq hz������ �
��.�@�m�d�v� ������ُЏ��� �*�<�i�`�r����� ��՟̟ޟ���&� 8�e�\�n�������ѯ ȯگ����"�4�a� X�j�������ͿĿֿ �����0�]�T�f� �ϊϜ����������� ��,�Y�P�bߏ߆� ���߼��������� (�U�L�^������ �������� ��$�Q� H�Z���~��������� ������ MDV �z������ �
I@Rv �������/ /E/</N/{/r/�/�/ �/�/�/�/�/??A? 8?J?w?n?�?�?�?�? �?�?�?�?O=O4OFO sOjO|O�O�O�O�O�O �O�O_9_0_B_o_f_ x_�_�_�_�_�_�_�_ o5o,o>okoboto�o �o�o�o�o�o�o1 (:g^p��� ���� �-�$�6� c�Z�l�������ϏƏ ؏���)� �2�_�V� h�������˟ԟ� ��%��.�[�R�d��� ����ǯ��Я���!� �*�W�N�`������� ÿ��̿޿���&� S�J�\ωπϒϿ϶� ��������"�O�F� X߅�|ߎ߻߲����� �����K�B�T�� x����������� ��G�>�P�}�t��� ���������� C:Lyp��� ���	 ?6 Hul~���� �/�/;/2/D/q/ h/z/�/�/�/�/�/? �/
?7?.?@?m?d?v? �?�?�?�?�?�?�?O 3O*O<OiO`OrO�O�O��O�O�F  �H551�C�A2��FR782�G50��EJ614�EAT�UPV545X6��EVCAM�ECU�IFW28[VNR�EV52NVR63�WSCH�ELIC�~VDOCV�VCS]UV869W0*V�EIOCW4VR{69NVESET7WvMWJ7MWR68�F�MASK�EPRXuYgX7�FOCOh�37XV`X3VfJ�6X53�VH�hL{CH>fOPLG7W�0nfMHCR?fS��gMAT~VMCS�6X0g55*VMD�SW#wagOPagM�PRbf�P�h0VPCMfW5iw`*V�`��g51BW51�x0nBVPRSg69Vf�FRDZVFREQnVMCN�F93V�SNBA�W�gSH�LB�M)��Px2�VHTC6VTMI�LX�VTPA�VT7PTX[�EL�v�`��W8WP�FJ95�rVTUTbfUEV�fUEC>fUFR�ZVVCC��O�fV�IPf�CSC��C�SG~V�PI�EWE�B6VHTT6VR6��X��3P>�CGU�I�G=�IPGS��RmCf�DGagH7�w��`W51�X6nh0HrVK�nh5NV�PJxj�x6rWL)�J7!�;R7�gS50W̘wJ64�VR55nf��rV�P�w76h7��FS�Z4��5ɧRm6�gR9٘79zh�4rV��VfWN	wR�8!wR76BW76�VfD06*VFL�R�TS�CRDfC;RXbfCLIRxAW�CMS�V��6VSTuYf�6!wCTO6V��P�W7�W�P�NN��VfORS�f/`VwFCB�VFCF�w�CH6VFCRfF[CI��FC�gJ��Z�gM�gPG�M�xwR58*VNETfV�NOM�VCp�VOP�a�SEND?fAP�>�PLU�f�P��7��VCPR�wL�S��C�Y67VfETaS�Ǡ��Pr�CP~V�TEq�S6]�TO�A.vTRA>fINv�wIHY�IPNf� �H������%�7�I� [�m��������� �����!�3�E�W�i� {��������������� /ASew� ������ +=Oas��� ����//'/9/ K/]/o/�/�/�/�/�/ �/�/�/?#?5?G?Y? k?}?�?�?�?�?�?�? �?OO1OCOUOgOyO �O�O�O�O�O�O�O	_ _-_?_Q_c_u_�_�_ �_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o �o�o�o%7I [m����� ���!�3�E�W�i� {�������ÏՏ��� ��/�A�S�e�w��� ������џ����� +�=�O�a�s������� ��ͯ߯���'�9� K�]�o���������ɿ ۿ����#�5�G�Yπk�}Ϗϡϳ������  H55������2��R78�2��50��J61�4��ATU��5�5�45/�6��VCA�M��CUIF/�2�8�NRE�52�n�R63�SCH���LIC��DOC�V��CSU�86�9/�0>�EIOC���4�R69n�EgSETO�m�J7m��R68�MASK^��PRXY��7��OCOo�3O��{��.�3��J6-�53��H�LCH��O�PLGO�0��MH�CR��Sm�MAT���MCSN�0~�5=5>�MDSW����;OP��MPR���к�0.�PCM��5`={�>�{��51^��51~0^�PRSvn�69��FRD~��FREQ�MCN���93.�SNBA����SHLBM�=����2.�HTC�N�TMIL��T{PA>�TPTX#EL�
{��8����J95��TUT���UEVn�UEC��UFR~�VCC�N,O��VIP�C;SC�CSG����I��WEBN�HTTN�R6���KЮ*�CG�+IG�+IP�GS:RC�DG���H7�+��51�N�6��0��k��5�n��J���6��L�=J7�;R7=�Ss50�l<J64�R55��[@��[�n�76~�7�S��4��5�KR6}�R9}<79��4�ګ@���WN��R8��R7�6^�76��D06�>�Fl\RTSC�RDn�CRX��CsLI]�CMS>�\�PN�STY�6��GCTON��>�7�̻О;NNNm��ORqS����.�FCB>�FCF�CHN�F�CRn�FCI.:F�C��J0��M��PuG�:M�R58>�wNET��NOM>�� �OP�kSEN�D��AP�*PLU�n��nL7�CPR��L]+S|lC�67��ETS~{�\+ඞCP��TE�[S�6-KTOA��TRmA��IN�IH}IPN���Տ��� ��/�A�S�e�w��� ������џ����� +�=�O�a�s������� ��ͯ߯���'�9� K�]�o���������ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ������� ����1�C�U�g�y� �ߝ߯���������	� �-�?�Q�c�u��� �����������)� ;�M�_�q��������� ������%7I [m����� ��!3EWi {������� ////A/S/e/w/�/ �/�/�/�/�/�/?? +?=?O?a?s?�?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O �O�O�O_#_5_G_Y_ k_}_�_�_�_�_�_�_ �_oo1oCoUogoyo �o�o�o�o�o�o�o	 -?Qcu�� �������)� ;�M�_�q��������� ˏݏ���%�7�I� [�m��������ǟٟ ����!�3�E�W�i� {�������ïկ��� ��/�A�S�e�w��� ������ѿ����� +�=�O�a�sυϗϩ���������S�TD��LANG����(�:�L�^� p߂ߔߦ߸�������  ��$�6�H�Z�l�~� �������������  �2�D�V�h�z����� ����������
. @Rdv���� ���*<N�`r���RB=T�OPTN�� �//%/7/I/[/m/ /�/�/�/�/�/�/�/�?!?3?DPN �Q?c?u?�?�?�?�? �?�?�?OO)O;OMO _OqO�O�O�O�O�O�O �O__%_7_I_[_m_ _�_�_�_�_���_ �_	oo-o?oQocouo �o�o�o�o�o�o�o );M_q�� �������%� 7�I�[�m�������� Ǐُ����!�3�E� W�i�{�������ß՟ �����/�A�S�e� w���������ѯ��� ��+�=�O�a�s��� ������Ϳ߿��� '�9�K�]�oρϓϥ� �����������#�5� G�Y�k�}ߏߡ߳��� ��������1�C�U� g�y���������� ��	��-�?�Q�c�u� �������������� );M_q�� �����% 7I[m��� ����/!/3/E/ W/i/{/�/�/�/�/�/ �/�/??/?A?S?e? w?�?�?�?�?�?�?�?@OO+O=OOOaH�aO�O�O�O�O�O�J9�9�E�$FEAT�_ADD ?	����
QP  	�H_-_?_ Q_c_u_�_�_�_�_�_ �_�_oo)o;oMo_o qo�o�o�o�o�o�o�o %7I[m �������� !�3�E�W�i�{����� ��ÏՏ�����/� A�S�e�w��������� џ�����+�=�O� a�s���������ͯ߯ ���'�9�K�]�o� ��������ɿۿ��� �#�5�G�Y�k�}Ϗ� �ϳ����������� 1�C�U�g�yߋߝ߯� ��������	��-�?� Q�c�u������� ������)�;�M�_� q��������������� %7I[m ��������DDEMO �
Y?   �HD :Lyp���� ���//?/6/H/ u/l/~/�/�/�/�/�/ �/??;?2?D?q?h? z?�?�?�?�?�?�? O 
O7O.O@OmOdOvO�O �O�O�O�O�O�O_3_ *_<_i_`_r_�_�_�_ �_�_�_�_o/o&o8o eo\ono�o�o�o�o�o �o�o�o+"4aX j������� �'��0�]�T�f��� ����ɏ��ҏ���#� �,�Y�P�b������� ş��Ο����(� U�L�^����������� ʯ����$�Q�H� Z���~�������ƿ� ��� �M�D�Vσ� zόϹϰ�������� 
��I�@�R��v߈� �߬߾�������� E�<�N�{�r���� ���������A�8� J�w�n����������� ����=4Fs j|����� �90Bofx �������/ 5/,/>/k/b/t/�/�/ �/�/�/�/�/?1?(? :?g?^?p?�?�?�?�? �?�?�? O-O$O6OcO ZOlO�O�O�O�O�O�O �O�O)_ _2___V_h_ �_�_�_�_�_�_�_�_ %oo.o[oRodo�o�o �o�o�o�o�o�o! *WN`���� ������&�S� J�\������������ ڏ���"�O�F�X� ��|�������ߟ֟� ���K�B�T���x� ������ۯү��� �G�>�P�}�t����� ��׿ο����C� :�L�y�pςϜϦ��� ����	� ��?�6�H� u�l�~ߘߢ������� ����;�2�D�q�h� z������������ 
�7�.�@�m�d�v��� ������������3 *<i`r��� ����/&8 e\n����� ���+/"/4/a/X/ j/�/�/�/�/�/�/�/ �/'??0?]?T?f?�? �?�?�?�?�?�?�?#O O,OYOPObO|O�O�O �O�O�O�O�O__(_ U_L_^_x_�_�_�_�_ �_�_�_oo$oQoHo Zoto~o�o�o�o�o�o �o MDVp z������� 
��I�@�R�l�v��� ����ُЏ���� E�<�N�h�r������� ՟̟ޟ���A�8� J�d�n�������ѯȯ گ����=�4�F�`� j�������ͿĿֿ� ���9�0�B�\�fϓ� �Ϝ������������ 5�,�>�X�bߏ߆ߘ� �߼��������1�(� :�T�^������� ������ �-�$�6�P� Z���~����������� ����) 2LV� z������� %.HRv� ������!// */D/N/{/r/�/�/�/ �/�/�/�/??&?@? J?w?n?�?�?�?�?�? �?�?OO"O<OFOsO jO|O�O�O�O�O�O�O ___8_B_o_f_x_ �_�_�_�_�_�_oo o4o>okoboto�o�o �o�o�o�o0 :g^p���� ��	� ��,�6�c� Z�l�������ϏƏ؏����(�   �>�P�b�t������� ��Ο�����(�:� L�^�p���������ʯ ܯ� ��$�6�H�Z� l�~�������ƿؿ� ��� �2�D�V�h�z� �Ϟϰ���������
� �.�@�R�d�v߈ߚ� �߾���������*� <�N�`�r����� ��������&�8�J� \�n������������� ����"4FXj |������� 0BTfx� ������// ,/>/P/b/t/�/�/�/ �/�/�/�/??(?:? L?^?p?�?�?�?�?�? �?�? OO$O6OHOZO lO~O�O�O�O�O�O�O �O_ _2_D_V_h_z_ �_�_�_�_�_�_�_
o o.o@oRodovo�o�o �o�o�o�o�o* <N`r���� �����&�8�J� \�n���������ȏڏ ����"�4�F�X�j� |�������ğ֟��� ��0�B�T�f�x��� ������ү����� ,�>�P�b�t������� ��ο����(�:� L�^�pςϔϦϸ��� ���� ��$�6�H�Z� l�~ߐߢߴ������� ��� �2�D�V�h�z� ������������
� �.�@�R�d�v����� ����������* <N`r��������&  '!BTf x������� //,/>/P/b/t/�/ �/�/�/�/�/�/?? (?:?L?^?p?�?�?�? �?�?�?�? OO$O6O HOZOlO~O�O�O�O�O �O�O�O_ _2_D_V_ h_z_�_�_�_�_�_�_ �_
oo.o@oRodovo �o�o�o�o�o�o�o *<N`r�� �������&� 8�J�\�n��������� ȏڏ����"�4�F� X�j�|�������ğ֟ �����0�B�T�f� x���������ү��� ��,�>�P�b�t��� ������ο���� (�:�L�^�pςϔϦ� �������� ��$�6� H�Z�l�~ߐߢߴ��� ������� �2�D�V� h�z���������� ��
��.�@�R�d�v� �������������� *<N`r�� �����& 8J\n���� ����/"/4/F/ X/j/|/�/�/�/�/�/ �/�/??0?B?T?f? x?�?�?�?�?�?�?�? OO,O>OPObOtO�O �O�O�O�O�O�O__ (_:_L_^_p_�_�_�_ �_�_�_�_ oo$o6o HoZolo~o�o�o�o�o �o�o�o 2DV hz������ �
��.�@�R�d�v� ��������Џ��� �*�<�N�`�r����� ����̟ޟ���&� 8�J�\�n��������� ȯگ����"�4�F� X�j�|�������Ŀֿ �����0�B�T�f� xϊϜϮ��������� ��,�>�P�b�t߆� �ߪ߼��������� (�:�L�^�p���� �������� ��$�6� H�Z�l�~��������� ������ 2DV hz������P�
,0# FXj|���� ���//0/B/T/ f/x/�/�/�/�/�/�/ �/??,?>?P?b?t? �?�?�?�?�?�?�?O O(O:OLO^OpO�O�O �O�O�O�O�O __$_ 6_H_Z_l_~_�_�_�_ �_�_�_�_o o2oDo Vohozo�o�o�o�o�o �o�o
.@Rd v������� ��*�<�N�`�r��� ������̏ޏ���� &�8�J�\�n������� ��ȟڟ����"�4� F�X�j�|�������į ֯�����0�B�T� f�x���������ҿ� ����,�>�P�b�t� �ϘϪϼ�������� �(�:�L�^�p߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v������� *<N`r� ������// &/8/J/\/n/�/�/�/ �/�/�/�/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $ 6HZl~��� ����� �2�D� V�h�z�������ԏ����
��.��$F�EAT_DEMO�IN  3���^��4�F�IND�EXS�b��F�I�LECOMP ߄������a�A���SETU�P2 ���~���  N ɑ���_AP2BCK� 1���  #�)/����%�0�4����[�1�򟇯 ���:����p���� )�;�ʯ_����$� ��H�ݿ�~�Ϣ�7� ƿD�m����� ϵ��� V���z��!߰�E��� i�{�
ߟ�.���R��� �߈���A�S���w� ���<���`���� ��+���O���\���� ��8�����n���' 9��]����"� F�j��5� Yk����T �x//�C/�g/ �t/�/,/�/P/�/�/ �/?�/??Q?�/u?? �?�?:?�?^?�?�? O�)O��אP۟ 2~�*.SPB0O�{O %FRH:�\PLUGIN\�eO1��0�O�O�5�*.VR�O�O�0* �O(_�2-_Q_�H�PCY_�_�0FR#6:mR_�Y=_�_�KTr��_o�U�P�_@2iU��_Xo�6d@F�O��o�1	�Swa'o�h8Eo�oikSTM�o �R�P�a&o:y�o^ikH�o� wq.@8��nfGIF���"u���Y�k�nfJPGq���"u��6�H�ݏ��FJS����0���S _ˎ
J�avaScriptJ�u�CS���!v���>�̍Casc�ading St�yle Shee�tsΟ�0
ARGNAME.DT����<%p\�ȟ҇��R����DISP*��>=���M��_���֯��CLL�B.ZI󯮯�`:�\�\�oZ�1�C?ollaboZ��
PANEL1�oി;���T�҇iP�endant POanel޿�8	������ɸ(�S�����ϛ�2����Ǹ��\�nπϒ� �2'�@�K�@.�[���ߘߛ�3�� ��Ǹ��d�v߈ߚ� �3/�H�K�6�c�����4����Ǹ��l�~��� �47�P�K��>�k�����)
T�PEINS.XML����:\��t����Custom T?oolbar�����PASSWORD<?��>FRS˱C�Passwo�rd Config��?�Z�O %�I[�� �D�h���3/ �W/�P/�//�/@/ �/�/v/?�//?A?�/ e?�/�??*?�?N?�? r?�?O�?=O�?aOsO O�O&O�O�O\O�O�O _�O�OK_�Oo_�Oh_ �_4_�_X_�_�_�_#o �_GoYo�_}oo�o0o Bo�ofo�o�o�o1�o U�oy��>� �t	��-���c� ��������L��p� ����;�ʏ_�q� � ��$���H�Z��~�� ���I�؟m������� 2�ǯV������!��� E�ԯ�{�
���.��� տd������/Ͼ�S� �wω�ϭ�<���`� r�ߖ�+ߺ�$�a��� ��ߩ߻�J���n�������$FILE�_DGBCK 1�������� < ��)
SUMMAR�Y.DG�U�MD�:M����Di�ag Summa�ry���CONSLOG��f�x�������� sole �lo���	TPA'CCN�l�%T������TP Acc?ountin3����FR6:IPKDMP.ZIP�����
�����Exception���y�MEMCHECCK����|�%��Memory D�ata���)�{�)�RIPE�pv��%�� Packet 9L2����\[�STAT��� %9St�atus�V	F�TP���/��'�mment T�BD*/�w��)�ETHERNE�o/\m/�/��E�thernB)�figura9��!?DCSVRF//�//?��  ve�rify all�2?��,�%DIFF'???�?3I8diff�?j7\� CHG01�?�?�?�9O��?aO����92/OO(O�O�?^O�pO�23�O�O�OA_� �Oh_�FVT�RNDIAG.LASm__0_�_��QO Ope�#D ��nostic���	l)VDEV�RDAT�_�_�_��_�Vis�QD�evice�_�[IMG�R$o6o�o2=adImagmo�[7UP`ESo�o?FRS:\R}���Update?s ListR����`FLEXEV�EN�/�o�o����q UIF Ev�E!E�{B�)�CRSENSPK�o����\��/� �CR_L�OR_P�EAKZ���PSRBWLD.CM�����=r��T&�PS�_ROBOWEL<K/�/:GIG�8���\��GigE��h��S�SAM���J�ߟ����/EmailcPa�����<<)ёHADOW۟��ҟg���Shadow Change���"C�'�RCMERR_�D�V�믮���CFG Er�rorg`t��� ���XcCMSGLIB�ʯܯq�0t�4��rpic�)�o�D)]�ZD��p˿Z�￪ZD���ad���Ό)v��T_�_RP��Կ���B�<��$ R�eport'�դ�7�IRDB�EPO�RF�X�j�|�%�iR�gs����N=t'�NOTI�/�����}߬Noti�fic�"��V��) ���<����p=���,�v�Y��� }����B���f��� ���1���U�g���� ���>�����t�	�� -?��c���( �L����; �4q �$�� Z�~/��I/� m///�/2/�/V/�/ �/�/!?�/E?W?�/{? 
?�?.?@?�?d?�?O �?/O�?SO�?LO�OO �O<O�O�OrO_�O+_ �O�Oa_�O�_�_&_�_ J_�_n_�_o�_9o�_ ]ooo�_�o"o�oFoXo �o|o#�oG�ok �od�0�T�� ���C���y�� ����>�ӏb������� -���Q���u������ :�ϟ^�p����)�;� ʟ_���|���H� ݯl�����7�Ư[� ����� ���ǿV�� z�Ϟ��E�Կi��� �ϟ�.���R���vψ������$FILE�_FRSPRT � �������7�MDONLY 1�K�~�� 
 ��� ���ϲ��Ͽ��߱�� ��0�B���f��ߊ�� +���O��������� >���K�t����'��� ��]�����(��L ��p��5�Y � �$�HZ� ~��C�g� /�2/�V/�c/�/~5�VISBCKi�|S�x�*.VD�/|�/K FR:\� �ION\DATA�\�/F"K Vi�sion VD file	?/Q?c? y/�?q/�?:?�?�?p? O�?)O;O�?_O�?�O O$O�OHO�O�O�O_ �O7_�OH_m_�O�_ _ �_�_V_�_z_o�_�_ Eo�_io{o6o�o.o�o Ro�o�o�o�oAS �ow�*<�1��LUI_CONF�IG �K�|�!�{ $ �sn�{K�3�E�W�i�{������|x�ŏ׏ �������@�R�d� v��������П��� ���*�<�N�`�r��� �����̯ޯ���� &�8�J�\�n������ ��ȿڿ�����"�4� F�X�j�|�Ϡϲ��� �����ϑ��0�B�T� f�x�ߜ߮������� {����,�>�P�b��� ���������w�� �(�:�L�^������ ��������s� $ 6HZ��~��� ��o� 2D V�z����� k�
//./@/�Q/ v/�/�/�/�/U/�/�/ ??*?<?�/`?r?�? �?�?�?Q?�?�?OO &O8O�?\OnO�O�O�O �OMO�O�O�O_"_4_ �OX_j_|_�_�_�_I_ �_�_�_oo0o�_To foxo�o�o3o�o�o�o �o�o>Pbt ��/����� ��:�L�^�p����� +���ʏ܏� ���� 6�H�Z�l�~���'����Ɵ؟������R�obot Spe?ed 10%�I��[�m������  �x�����$FL�UI_DATA �����ա���ǤRESULT 3�ե��� �T��/wizard�/guided/�steps/Expert��5�G�Y� k�}�������ſ׿�����Conti�nue with{ G�ance�� 2�D�V�h�zόϞϰϰ�������� ���-��ե�0 a����A�ա�	�ps�ςߔߦ߸��� ���� ��$�6�H�� ��o��������� �����#�5�G���ᢠ��G�)ߋ�M�]�c�llb�Sele?ctWorkP��� ��'9K]o�����Ligh�twe� ��pie����1�CUgy��� a�y����&]��rip ��Too�lNum/NewFram�;/M/_/ q/�/�/�/�/�/�/�/�0x0�/?-? ??Q?c?u?�?�?�?�?8�?�?�?  �����3OM�]�!imeUS/DST�? �O�O�O�O�O�O�O_�_+_=_ �Enabl*/q_�_�_�_�_ �_�_�_oo%o7oIo���!O�o�oWOiF24tO�o�o�o !3EWi{�L_ ^_������/� A�S�e�w�����Zolo�~o��R���ditor��-�?�Q�c�u����������ϟ��� �Touch Pa�nel � (recommen�)�4�F�X�j�|��������į֯�ب�����ɏ+�=����accesp߀������� ȿڿ����"�4�O��Conn�� t?o Netw��w� �ϛϭϿ���������+�=߬�_�?�!����!U��Int�roductionF��������#�5� G�Y�k�}����|Ь� ����������*�<� N�`�r��������O�pߒ�����4��c�llb�Load�SettingN?otHW_l�"W���BTfx���������.0 �'9K] o��������	O������-/��8���!CenterMan��/�/�/�/ �/�/??(?:?�^? p?�?�?�?�?�?�?�?  OO$O6O�//{O�O�5Q/c/u(�0 �O�O_ _2_D_V_h_�z_�_��EOAT� w/o par �O�_�_�_�_oo0o@BoTofoxo�o��UO���o�o��+�O&�D�/DistanceWf�2DVhz ������Q?
� �.�@�R�d�v����� ����Џ�MO_OqO'���&�oz'Off ꏄ�������̟ޟ�`��&�8�S�1;� a�s���������ͯ߯@���'�9��
��"��oy���%M�_� ��ֿ�����0�B� T�f�xϊ�I�2�ϵ� ���������!�3�E�@W�i�{ߍ�L��k����?..��/�@Sp�eedLimit/Max��4�F� X�j�|���������Z	1�p���0� B�T�f�x���������0��������Dz�#�A,��guide}d�afety�� u������� )�[�N`r �������/ /&/8/g����oW/�/|CURegioſ �/�/�/�/?"?4?F?�X?j?|?�\UTC�+01 ~ �23 �?�?�?�?�?OO+O@=OOOaOsO�O��M"�}���/i/�O����/	qimezone5�O _2_D_V_h_�z_�_�_�_�_�_��<�(�3:00) A�m��rdam, ?Berlinb`�Rome, St�ockhol`Vienna�_@oRo dovo�o�o�o�o�o�OM!�ѾүO�O#�/�Oe24�oq�� �������%� <I�[�m�������� Ǐُ����!�3�J/�x���#EWv/?curren"�̟ ޟ���&�8�J�\��n�����17-JUL-24 1�P9 ����ί��� �(�:�L�^�p�����A��[���Ͽ�� ����Year���0� B�T�f�xϊϜϮ�������20^�� &�8�J�\�n߀ߒߤ߀���������a�����跿!��Month��s��� �����������'���7/�U�g�y��� ������������	-���� �m��9A𧻓Day2� ���1CUgy��1C��� ���//'/9/K/ ]/o/�/@R	_�/8ۿ���Hou�? +?=?O?a?s?�?�?�?�?�?�1�?�?O"O 4OFOXOjO|O�O�O�O�O�O�/S�/_���"�/S�inute �Op_�_�_�_�_�_�_ �_ oo$o;�9+oQo couo�o�o�o�o�o�o@�o)�OR		_�i��.=Ucllb���SetSpeedLimit/�wVal.������*�<�N�`�r���250.0����� ��Џ����*�<��N�`�r���A{uCz  _�����rMod^_�&�8�J� \�n���������ȯ���Do not �Use (Rec_ommen��)ӯ �"�4�F�X�j�|���p����Ŀ־ 8p�"8pϟ]�-\)��/Load�pt�ingNotHW?_lightֿs� �ϗϩϻ�������� �ԯZ=�O�a�s߅� �ߩ߻��������� '�8q걚� �"�t���abSummar����������� (�:�L�^�p�/ߔ��� �������� $6 HZl~=�O���5T#��file2�/cyclepowerKTm�$ 6HZl~���<��6HOT�� 	//-/?/Q/c/u/�/`�/�/�/�/�!����?-\9�/ToolP��/d?v?�? �?�?�?�?�?�?OO ��<ONO`OrO�O�O�O �O�O�O�O__&_��/A_k_�� 5?�{(_ �_�_�_�_oo&o8o Jo\ono-O�o�o�o�o �o�o�o"4FX�j)_;_M_�����_/����%�7�I� [�m��������Ǐ�o ����!�3�E�W�i� {�������ß������(�/Con�figurati�onCompleti�{�������ï կ�����܏A�S� e�w���������ѿ�����ח���?��iχ�XIntroducM�$ϵ����� �����!�3�E�W�i� (��ߟ߱��������� ��/�A�S�e�w���Hϒ��.<guid�ed�tNetMethodx���,� >�P�b�t���������~�Not cE�e����/AS�ew����~�  ���ŭ�= Oas����� ��//��9/K/]/ o/�/�/�/�/�/�/�/�/?�� �;? e?'�?�?�?�?�?�? �?
OO.O@OROdO#/ �O�O�O�O�O�O�O_ _*_<_N_`_?1?C? U?�_y?�_�_oo&o 8oJo\ono�o�o�o�o uO�o�o�o"4F Xj|�����_ �_�_	��_0�B�T�f� x���������ҏ��� ��o,�>�P�b�t��� ������Ο����� ���[�������� ��ʯܯ� ��$�6� H�Z��k�������ƿ ؿ���� �2�D�Vπh�'���K�������n�etwork��AutoDHCPm�  ��$�6�H�Z�l�~� �ߢߴ�s��������  �2�D�V�h�z�������Ϝ�����&�����/robotip��\�n������� ������������4 FXj|���� ���u�����U��%%�7�status��� ��	//-/?/Q/c/>"ailedg/�/ �/�/�/�/�/�/?"? 4?F?X?);�?�?zu�ycllb�� j?�?OO&O8OJO\O nO�O�O�O�O!�O�O �O_"_4_F_X_j_|_�_�_�_�Z?�?�_�ow�ygripper�?AoSoeowo �o�o�o�o�o�o�o �O+=Oas�� �������_�_ �_0�Z�x��������� ɏۏ����#�5�G� Y�}�������şן �����1�C�U�p� ^�8�J���n� y���settingsp2e�����0�B� T�f�x�������m�ҿ �����,�>�P�b� tφϘϪ���'�������sկp2/name��S�e�w߉ߛ߀�߿��������ƱROBOT�5�G� Y�k�}�������� �����|?����R�l��&!o�ToolN�um/Fr?�Us Aߧ���������`%7I[Ʊ1_ �������@'9K]��
!� ;���;��n)q���?Active��b �/#/5/G/Y/k/}/x�/�/`
0xf�$ �/�/�/??*?<?N?@`?r?�?�?�?�:�������?��ܠM�acro��s/New/B5oROdOvO�O��O�O�O�O�O�O_�0x0_/_A_S_ e_w_�_�_�_�_�_�_��_o�6'��?CoUo��,O+K/BOpen ���o�o�o�o�o %7I_r�� ������!�3��E�W�n�:o��^k-|moooClos�� ����1�C�U�g�y�����\�ԟ��� 
��.�@�R�d�v�������k�}����[n9��/�Set/B�� D�V�h�z�������¿0Կ���YYeAO*� <�N�`�rτϖϨϺϠ������߼ �!A���+o�G�ah�>'�ethodߙ� �߽���������)��;�M�'Dire�ct entry� of EOAT dataW��� ����������%�7� I�߼!�"�4ߖ�\m�$i�'�traig�htOffset Z���(:L^�p����"��  ����%7 I[m��b��v����\m%������%%X�G/Y/k/}/�/��/�/�/�/�/�/�.00�/)?;?M?_? q?�?�?�?�?�?�?�?Oů� �AO//'+YO�O�O�O�O �O�O__+_=_O_? s_�_�_�_�_�_�_�_ oo'o9oKo
OO.O0�oROdOvOtZVo�o %7I[m ��b_����� !�3�E�W�i�{����� ^opo�o䏦o)�o���Rotation!�W��G�Y�k�}��� ����şן韨�� 1�C�U�g�y������� ��ӯ�����ȏڏ<����"�nP������ ��ѿ�����+�=� ���sυϗϩϻ��� ������'�9�K�
���.���R�d�v�nR R�����%�7�I�[� m���P�b������� ���!�3�E�W�i�{������^�p߂����k"�����tp3Zdi?r/Tp3z��< N`r����� ����&8J\ n�������@��������C/�`+	���Measure�ment/Straigh�o�/�/�/ �/�/�/??'?9?� 
o?�?�?�?�?�?�? �?�?O#O5OGO//p*/�ON/`//We�!�Nums/New�CsNO�O�O_#_5_�G_Y_k_}_�_N=0xc?�_�_�_�_o o 2oDoVohozo�o�ob@AaO�iO�o��.�O��LTool�CUse�oDVhz��`����Q:1� �+�=�O�a�s�����@����͏ߏ�a
�o�wD�o1��o�LPart*������ş ן�����1�C��2G�m��������ǯ ٯ����!�3�E��"rI#�����(Y��Gs/G���CJ���� 
��.�@�R�d�vψ� ��]?���������� *�<�N�`�r߄ߖ�YO�kO}O����)����P�ayload1CmԿ:�L�^�p�������������E�OAT w/o p{���!�3�E�W�i� {������������������o7���x� ����������0B�10 ��j|����� ��//0/B/��?	�A �߃/��W�2 '��/�/??(?:?L?�^?p?�?�?���ith��?�?�?�?O O1OCOUOgOyO�O�� \/�O�OP&�/�)�Advanced �O4_F_X_j_|_�_�_�_�_�_�_��0x ]o$o6oHoZolo~o��o�o�o�o�o�o�@ �O�O	3Q�%�O�!�Mass/Centergq�o��� ������)�;� ��_�q���������ˏ ݏ���%�7�N/`��|�>�/bsss B�ߟ���'�9�K� ]�o���@�R���ɯۯ ����#�5�G�Y�k��}���N�`�r�Կ��,����!GPcmr��X ��6�H�Z�l�~ϐϢ� �����ϗ���� �2� D�V�h�zߌߞ߰��� ���ߥ���ɿ+�����sY�ߊ����� ��������,����� b�t������������� ��(:����0A�S�e�sZ>� �&8J\n �?�Q������ /"/4/F/X/j/|/�/ M_q�/��.�� �1��$�3?E?W?i?{? �?�?�?�?�?��O O/OAOSOeOwO�O�O �O�O�O�O�/�/�/(_�/�/?rtx�_�_ �_�_�_�_�_oo)o �?�?_oqo�o�o�o�o �o�o�o%7�O�__|>_P_b_rt �����#�5�G� Y�k�}�<oNo��ŏ׏ �����1�C�U�g� y���J\nП��|�TCPVerif�y/
�Method��.�@�R�d�v����������Я��Di�rect Entry߯�"�4�F�X� j�|�������Ŀֿ��A������!Ϗz'��fy"?|ώϠϲ� ����������0ߛ� T�f�xߊߜ߮����� ������,ϻ�0q�3�E�W�fyv_�� ������*�<�N�`� r���Cߨ��������� &8J\n��?�m�c������fy�$6HZl~ ��������/  /2/D/V/h/z/�/�/ �/�/�/���?���fyW�/y?�? �?�?�?�?�?�?	OO -O�QOcOuO�O�O�O �O�O�O�O__)_�/��/?n_0?B?T?yP 2_�_�_�_oo'o9o Ko]ooo�o@O�o�o�o �o�o�o#5GY k}<_N_`_��_�_�_yR�!�3�E�W� i�{�������ÏՏ�o ����/�A�S�e�w� ��������џ������}*��fyMeanڟx����������ү�����َ*?�+�X�j�|����� ��Ŀֿ�����ݟ �M��m��z)=�O�a�ax.�������� �%�7�I�[�m�,�>� �ߵ����������!� 3�E�W�i�{�:�|�^�����{"�ϣ�Int�roductio f��)�;�M�_�q��� ��������������  2DVhz� ������������r#��fil�e2/cycle�pow��done �m����� ��/!/��E/W/i/ {/�/�/�/�/�/�/�/??,;��G?q?��r,��crsgd�etail��Se�lectCate�gory/list,?�?�?�? OO$O�6OHOZOlOیAl�loc�0d by? KAREL{O�O �O�O�O�O__0_B_PT_f_x_�����Q�w?Y?�_�|/�?��_force/F�Q?Limit1�?o .o@oRodovo�o�o�o|�oَ--- �O �o
.@Rdv ������T�R�_@�_��_�_�_`2o p���������ʏ܏�  ���o�o#�Z�l�~� ������Ɵ؟����  ��!��e�'�9�K�t3_�į֯���� �0�B�T�f�%�7�w� ����ҿ�����,� >�P�b�t�3�u�W���{�����t4���*� <�N�`�r߄ߖߨߺ� y�������&�8�J� \�n�������ϐ�ϫ��+6����p�ayload�4P�K�No/check��x�����������`������  �O EWi{���� ���������^ �71�C�ldc�hg/P�Ena�bleSignal�����/"/ 4/F/X/j/�O;�/�/ �/�/�/�/??0?B?PT?f?%�Pb�Po�Q�?!����spd�lmt/S�2Clamp��O-O?O QOcOuO�O�O�O�O���Њ/�O__%_7_ I_[_m__�_�_�_�_ ��?�?o�78�?�5tatus/SGb�Safety�1 
Oqo�o�o�o�o�o�o �o~/�OI[m ������� ��_�_�_<�f�(o:oLol2`oŏ׏��� ��1�C�U�g�&8 ������ӟ���	�� -�?�Q�c�"�4�F���0��|�����l3��� +�=�O�a�s������� ��z������'�9� K�]�oρϓϥϷ�v���������Я���l4�m�ߑߣߵ���`��������E-�@ ۿ@�R�d�v���� ��������������@��]��1�C߱5\� ��������	-? Qcο4���� ��);M_@�0�B����19}����usDigitalYo/!/3/E/W/ i/{/�/�/�/p��/ �/??/?A?S?e?w? �?�?�?�?~c�� �?O�����iO{O �O�O�O�O�O�O�O_ �/�/A_S_e_w_�_�_ �_�_�_�_�_o�?�? �?4o^o O2ODO��o �o�o�o'9K ]_._����� ���#�5�G�Y�o *o<oNo��ro�o�oW� ��1�C�U�g�y��� ����n����	�� -�?�Q�c�u������� ��|������ď֏� ��_�q���������˿ ݿ����ҟ7�I�[� m�ϑϣϵ������� ���ί��T��(�:��6U��������� ��&�8�J�\��-� ������������� "�4�F�X��)�;߅���q�)u߇�ats�ts/A��Checkf�'9K�]o���d�DISABLE � ��,>Pb�t����k�d0����/�+����?TimeLm��X/ j/|/�/�/�/�/�/�/ �/��?B?T?f?x? �?�?�?�?�?�?�?O �	/�MOg�5///InputA$�߲O �O�O�O�O__0_B_<T_k�-- z�_ �_�_�_�_�_�_oo )o;oMo_ov�0OBO�o�j�0qO�OWarning�O%7 I[m��f�x�s��)����(� :�L�^�p�������eo��pˁ�o�o�e�*��o�frsm��4�Enable��T�f� x���������ҟ��� ??�>�P�b�t��� ������ί���O���I�g�3�+�PrgRun�o���� ̿޿���&�8�J� ��[ϒϤ϶����� �����"�4�F�X�ooY�;���cJ1m����Pause����� "�4�F�X�j�|��� _�q���������0� B�T�f�x�������mߐߑ���eH%���c/�Introduction��K]o �������� ����5GYk}� ��������΁ ����C/aL!'CompletB� �/�/�/�/�/�/?? *?<?N?�?�?�? �?�?�?�?OO&O8O�JO��/-/wO�O�)|i/�dforce-F�AZO�O	__-_?_ Q_c_u_�_�_X?j?|? �_�_oo)o;oMo_o qo�o�o�ofO�O�O�o�^�/�O�J�BLim�it1/var1 �oQcu���� ����_�_)�;�M� _�q���������ˏݏ ���o�o�oF�,{2;����ğ֟� ����0�B���S� ��������ү���� �,�>�P��Q�3���W�i�{�t3����� �*�<�N�`�rτϖ� U�g���������&� 8�J�\�n߀ߒߤ�c�������߫���Ͽt4 �H�Z�l�~���� ������ϻ���2�D� V�h�z����������������������=��.|��JEscap4s 7��������� 0B��x� ������// ,/>/P/!3�/��+a�JSummary�O�/�/?"?4? F?X?j?|?�?�?_q �?�?�?OO0OBOTO fOxO�O�O[/�//�O���(�/�Comp �/=_O_a_s_�_�_�_ �_�_�_�_�?�?'o9o Ko]ooo�o�o�o�o�o��o�o�O�O�O�OD���-	_�payl�oad/IntroPws�o���� ����+�=��_o s���������͏ߏ� ��'�9�K�
.䐟�5]o|Sel7ect�tNo7�� ��(�:�L�^�p��� ��S�e�ʯܯ� �� $�6�H�Z�l�~���O� a�s�����3��o|>�tWeigh�� H�Z�l�~ϐϢϴ��� ���ϩ��� �2�D�V� h�zߌߞ߰�������@����ɿ�=�[0��yqXYZ3ϕ�� ����������%�7� ���m���������� ������!3E��(�Py4Y�k�yqInertia�� ��#5GYk }�N�`����� //1/C/U/g/y/�/@�/\n��/Tu/�~Ýummary� :?L?^?p?�?�?�?�? �?�?�?��$O6OHO ZOlO~O�O�O�O�O�O@�O�/�/�//_M|,?o|Comp)?�_�_ �_�_�_�_�_	oo-o?nb�?Ovo�o�o �o�o�o�o�o*<<�1mers__�'_�KV+U_gUld�chg/IntroP�rA��	���-�?�Q�c�u����8gTooUogȍޏ�� ��&�8�J�\�n���~��  timeWi{ݟKV1��{�s?LimitX�:� L�^�p���������ʯܯ�7 ������ �2� D�V�h�z�������¿ Կ��O�ɟ+�����#�Y)��Ϡϲ��� ��������0��?� f�xߊߜ߮������� ����,�>����!�0��E�W�i�tZ}��� ����*�<�N�`�r� ��C�Uߺ������� &8J\n�� Q�c�u��IX6���!�Rot����;M _q������ ����/%/7/I/[/m/ /�/�/�/�/�/����?0?NS-��{S?ummary��? �?�?�?�?�?�?OO 'O9O�
/oO�O�O�O �O�O�O�O�O_#_5_ �/"??z_�}*M?�{Compt?�_�_�_ oo0oBoTofoxo�o IO[O�o�o�o�o ,>Pbt�E_W_�i_���+�_�Ts�pdlmt/IntroS��1�C� U�g�y���������ӏ �o�o	��-�?�Q�c� u���������ϟ០��&��Y2����Value/rw +��������Я��� ��*����`�r��� ������̿޿��π&�8���	��}ϗV7�I�[�mtClam�pEnabls�fl�_������,�>� P�b�t߆�E�W����� ������(�:�L�^�p��A�S�e�������5�ϯ�mtMaxSpeedt�0�B� T�f�x����������� �ߣ�,>Pb t�������� ����%C?��c�n3� }������� //1/��g/y/�/ �/�/�/�/�/�/	?? -?�r?�_F� �Ql�?�?�?OO(O`:OLO^OpO�O4C/ U/�O�O�O�O__&_ 8_J_\_n_�_??m?c?��_��?�tatus�b�_)o;oMo_o qo�o�o�o�o�o6/�O %7I[m ������_�_�_ �8�_feoz��� ����ԏ���
�� .��o�od�v������� ��П�����*�� +��o��?C�i�2i� ˯ݯ���%�7�I� [�m��>�P���ǿٿ ����!�3�E�W�i�@{�:�L�^��ς�)��^�4atstdA� ��#�5�G�Y�k�}ߏ� �߳��߄������� 1�C�U�g�y���� ������϶���_�� ��e�t��������� ������(���� ^p������ � $����i��(=��ʹ1c��� ��//1/C/U/g/ y/8J�/�/�/�/�/ 	??-???Q?c?u?4�FXz�?��L�rsm� @�?O1OCOUO gOyO�O�O�O�O�/�/ �/	__-_?_Q_c_u_ �_�_�_�_�_�?�?�? o.��?�7\�Oro�o �o�o�o�o�o�o &�O�O\n��� ������"��_ #oog��;o�8�ao ÏՏ�����/�A� S�e�w�6H����џ �����+�=�O�a�@s�2�D�V���z�'���O�/Select=C��gory~�� +�=�O�a�s���������Ϳ ������� �,�>�P�b�tφϘ� �ϼ�����˯����<�&�networ�k�settin�gsp2/ipadd��l�~ߐߢߴ߀��������� 
10.7� ?�D�V� h�z���������� ��
����	���a��>ᯣ&��������� ��0BTfѿ w�������,>Pbt���;�M����2��g�uided�NetDone|
// ./@/R/d/v/�/�/�/ �/}�/�/??*?<? N?`?r?�?�?�?�?�? ���O��5���Port�?\OnO�O �O�O�O�O�O�O�O_��GA 1 (CD38A)_R_d_ v_�_�_�_�_�_�_�_�oo�� ���B��O�?_o}�1O>��curit��o �o�o�o�o1C�Ug��?��L�ow (R-30�<i>i</i>B SL�@_��� ����1�C�U�g�^��o-ca3d����ooQo����os/methoZ��� )�;�M�_�q����������'V = n��Manual icß����+�=�O��a�s���������̗1073d��1Ï����%�ُ�bummar�oZ�l�~������� ƿؿ����͖)��/ >�P�b�tφϘϪϼ����������  eatu;a�?�;�e�8'���TesJO�� ����������,�>�8P�b�#� en-ϒ� ������������"��4�F�X�j�  tech'P3�Eߏ����� ���s�tp1 m�*<N`r�����ђope ����
.@R�dv����  age(/ߕ���	/�{f���Intro�U/g/y/�/�/�/��/�/�/�/	?'V800)�:?L?^?p?�? �?�?�?�?�?�? OO?  penV����]O{f%)/��/nameO�O�O�O�O��O__1_C_U_g^g�() �ROBOTg_�_�_�_�_�_ �_oo%o7oIo[oȞ� u�gOIO�oq�&<}O�Lipad� +=Oas����l�igh�1�92.168.150.2���� '�9�K�]�o���������u��o�o�o�w�9'�o�Lsub5��� ]�o���������ɟ۟�����59-1�_255.'�0� E�W�i�{�������ï�կ����z�m',�ӏ���Y��-��Drouter���ÿ տ�����/�A�S�c�0);
�{���� �ϼ���������(�p:�L�^�w�ady'��9�K���&$y��Lmace���&�8�J��\�n�����72�, �00:e���4:7d:bc:db������'� 9�K�]�o��������� {
  {ߍߟ�o��ߗB2E�Rd v�������<Addr %�2 DVhz���� ���
/y`������ ��U/);���/�/ �/�/�/??%?7?I?�[?@Quer�  �x/�?�?�?�?�? �? OO$O6OHOZOoSn=mi#/5/G/�O ��}/;���O__1_ C_U_g_y_�_�_�_xa �P���O�_�_o"o4o�FoXojo|o�o�o�o  ><imwO�O�O �ok&�`0BTf x�������� 4.�@�R�d� v���������Џ�� ��e�	�o-�W� ~�������Ɵ؟���@� �2�D�V��T0o� ��������ʯܯ� ���$�6�H�Z�  
[ 1�1�C���k&�#�O��NetTe�st/ipadd ]�����/�A�S�e��wωϛϭ� s)[/]�1x82���� ��	��-�?�Q�c�u� �ߙ߫��V�o�������k&&ſ׹linkstaGO�a�s�����������A�R-2�	Connected "� '�9�K�]�o������� �����������������D�!�׹url �������/ASg0WAR�N�http://�χ���� ��//)/;/M/�[A3-?�/�m װY/�/�/??/?A?�S?e?w?�?�?�<" DAq��?�?�?OO ,O>OPObOtO�O�O�O.�P000�s/�/ �O�Ok� _2_D_V_h_ z_�_�_�_�_�_�_�_�0 " _&o8o Jo\ono�o�o�o�o�o �o�o�os��O�OI _p�������� ��$�6�H��12:p�y��������� ӏ���	��-�?�Q� r�4��X��ϟ� ���)�;�M�_�q�x�������l?��� ί����(�:�L� ^�p�������e�ǿ�� 뿭��$�6�H�Z�l� ~ϐϢϴ����������\�� �2�D�V�h� zߌߞ߰��������� b�@��ѿ�E��l� ~�������������� �2�D�[�IS ic�v����������������*<N  vis=�%�7� �[����� ,>Pbt��[�id="����  //$/6/H/Z/l/~/��/�/  /cel gy��/�?&?8? J?\?n?�?�?�?�?�?x�?�?[�dius? O0OBOTOfOxO�O�O��O�O�O�O�O� dir�/�/�/A_?h_z_ �_�_�_�_�_�_�_
opo.o@o��loc__ ro�o�o�o�o�o�o�o�&8J  FAN�� _2_�V_� �����'�9�K��]�o������.00 �Ə؏���� �2� D�V�h�z������q�ew�����$F�MR2_GRP �1���� �C4  �B��	 �x1�C�.�F@ Y�y@�.�G�  ���Fg�fC�8R<��q�?�  �����.�6�X�Ѣ�8�75t��5��ߛ5`+�q�A�3  ���BH�o��%�@S331���-�S�d�.�@.�z�p� d�����ֿ������ 	�B�-�?�x�cϜ����_CFG ��TC�������
߬��NO �E169511��RM_CHKTYP  ��������ROMY�_MsIN_������u�J�X�SSB����� /��������߰��TP_DEF_O/W  ����ןIRCOM^����$GENOVRD�_DO����=�TYH���� dZ�dC�o_ENB/� C�RAVC������ �Q�H!�����ТI���PI\ٳI.��}������}����r�w��E� [��OU���� ��A��A�<ڒ����?�����|����C�  %���'9B���#D����ߤ�SMT����� ��Ч���$HOSTC��1�������� 5	�����	��e$Ugy ���C�����/�	anonymous/G/Y/k/ }/�/������// 1�$?6?H?Z?�~? �?�?�?�?�//-/O  O2ODOVO�/�/�/�/ �O�??�O�O
__._ q?R_d_v_�_�_�O�? O�_�_oo*omOO �O�O�_�o�O�o�o�o �oE_&8J\n �o�_�_����� AoSoeowoyj��o�� ����ď֏���� 0�S�A��x������� ��ҟ�'�9��M�>� ��b�t�����ۏ��ί ���'�(�k�L�^��p�����ן����18736��"�D� %�7�I�[�mϰ��ϣ� ��������.�@�!�3��E�W�i߬���SM
���ӷ5޿����� ����+�=��a�s� ��������������'�9��
�ENT� 1��	�  �P!ros p�cE�����!�192.168.�150.10��  !������������ &��Jn1�U ������4 �X-�Q�u �����0/�T/ /x/;/�/_/�/�/�/ �/�/?�/>??b?%? �?�?[?�??�?�?O��?(O�?�?^O!AQ�UICC��=O!%��2�OqG1�O�O'!
1���B �@�O�rF�O�OOOP_s@ROUTERR_._�K�O~ BPCJOG�_�}_!  ��^C�AMPRT�_�_!1���_�YRTk_o�/o�o !Sof�tware Op�erator P�anelmo!��G0 3�oT�NA�ME !c�!ROBCONT_�N�S_CFG 1��c� ��Auto-st�artedŴFTP �yq�߹� �������Y�4� F�X�j��{�!���ď ֏������Rdv W����n�����ß՟ ������/�A�d�� w���������ѯz߼� η��R�C���g�y� ������r�ӿ���	� ,�ƿ��Q�c�uχϙ� ��� ����&��Z� ;�M�_�q�4�.ߧ߹� ���� ���%�7�I� [�m����������� ����!�3�E��i� {���������V����� /A����� �������� ��=Oas��* ����//Xj |���/��/�/�/ �/�/�?#?5?G?Y? |/�/�?�?�?�?�?�? ,/>/P/Od?UO�/yO �O�O�O�O�?�O�O	_ _>O?_�Oc_u_�_�_�_3RI/&_ER�R �z�_�VP�DUSIZ  j3P^j@��T>�U?OLL ��_.@�  �I��` �6��UWRD �?@u-A�  �guest 3Vro�o�o�o�o�o.t�SCD_GROUoP 3�@| Dq�"IIFT~$P�A~OMP~ �~_SH~ED� ~$C~CO�M�PTTP_AU�TH 1�.k �<!iPend�an�g�~zF�!KAREL:*���}KC�#�5���VISION SET�`��j��������
��� @��)�K�M�_�\q�tCTR*`�.mB`Ζ�3Q
n��FF�F9E3��+DF�RS:DEFAU�LT�FAN�UC Web Server0ZߐΓ �tZold��g�y�����������TWR_CONFIG �u7�Q���Q�IDL_CPU_kPC�3QB�.@�3� A��_�M�IN$�	q >n��^�GNR_IO��Qb3P4h�HMI�_EDIT ��{
 ($fo�rlead	�0Z$7cu.� h���straig̿���regi  �ne����labe9lϵ�if��E�~�jump iD��޽kakujik�u�ϸ�	unde�f�������ݑ($ ��B�4q1�j�Uߎ�y� �ߝ����������0� �T�?�x�c�����2ROS2,1�49129630?1  069��/[����NPT_S_IM_DOi�s��NSTAL_SC�RNi� � �TPMODNTOL6��L�RTY�3�$�\���pENB6�	s��OLNK 1�.k�p��������� 2��MASTE�h���˒��SLA�VE �.kH �D��SRAMCA�CHEPb�qO_gCFG��	UO�����CMT_OPp�k�2j�YCL��
�_ASG 19����Q
 4W i{��������////A/<*N�UMc2i
�I�P��RTRY_�CN�2�_UP(� a����U �� F������̔�)��P0�?�.k ����F?X?j?|?�? �?;�5?�?�?�? OO $O�?HOZOlO~O�O�O 1O�O�O�O�O_ _�O �OV_h_z_�_�_�_?_ �_�_�_
oo.o�_Ro dovo�o�o�o;oMo�o �o*<�o`r ����I��� �&�8���n����� ����ȏW�����"� 4�F�Տj�|������� ğS�e�����0�B� T��x���������ү a�����,�>�P�߯ 񯆿������ο�o� ��(�:�L�^��� �Ϧϸ�����k�}�� $�6�H�Z�l��ϐߢ� ��������y�� �2� D�V�h���	����� ��������.�@�R� d�v������������ ������*<N`r ������ �&8J\n� !�����/� 4/F/X/j/|/�/(3�TIMER�#�!,��%�"_MEMBE�RS 2��%]�  $#5�"��),�'�/9� �RCA_ACC �3��%�!  � X�cZ ��[  -� 6�_� 6�n 6 ��!Q6	> -3�0a?S5 !"�<�34BUF001 �3�@;= ���u0  u0��*�4��4��3��0�2� �4@�4`�4�4���4��4��4��4���4�D�D��4���4��4��4��4���4�D�D��4���4��4��4��4���4�D�D��4���4��4��4��4a�Z]  ]a�zu@�^xaU��D��D��D��3�b$T:$TZ$TyT$TTbTbTb#T�c+Tc3Tc;TcpOP  OP��4U��4��4��4�D	�D�92�?�?�?�? OO*O<ONO`OrO�O��O�O�O�O�O�Kg{[�Q
�jP
_<_.Ud��:Q�Q BQGrpGrpGr$pGr ,p�QjQor3PorDt�Q �Q�_�_�_�33�_�U�  �S�p�R�p�R  �S�b�b�b���t#c��t3c   ;cB��KcB��[cB� �tkcB��t{c����c ����c���t�c���t �c��c��c`�t�c�t�C  �C 
�P�r
�r
�$r 
�,rIp+RIp3RIp;R Is8��RSas8�5�jS ysx�M��S�u& �t�s��p��s�p�34CF�G 3�@; 4��!�% < p�	��"34HIS�2ݧ@; �Q1 �2024-07-;18& �/l� ~�����#S0�ïկx���,X� C�!7O�Z�	��";V�� @�(@��r	�N�D�D�	�H@���	�X@��`8�f��p@�x
@��8��8���п���}C��1.�@� R�	��r �g�y����B �hğ�	�����U�ĘĠĨĵ�ĸĿ}�����5� ��Q�c�Q� ��sυ�����	��ϭ�p����	����`C� ���������	�� !�3���c�Q�cޘφӀ����	�����������3��������^� (�:�p����	�c��
;���2����+�=� 	������	���� ��K�9�o����P-��?�Q������� 
 2 �� ����������� 9 ��i �d��	�d�����'  C�����/ ��\n7ϒ���� �ߵ�������F/ |j/3�Eߠ/!��/�� �߱�?����B?�/ x?A�?/��,/�� OOP?>OPObO+��O �?a�s��?������:O ����pO^_�O9&��p Rdv�o�o�o�o� !�o,>P> �Lr�r$0r�@r �@r�pr�`r�r Pr��r��r��r ��r��r�r `r ��'�/'/�� ����,P��x(` �0`�8`��0��  �� �� �� ���/ T�f�x���������ҏ ����bq�?0�B�T� f�x���������ҟ�`_��O��0�B�T� f�x��������bq�_ �����0�B�T�f��x������ CI_C�FG 3�xk �H
Cycle� Time��Busy�I�dl����minz���Up�ƾ��Read���Dow���� �����Count>��	Num ���Ñ��]�� 5�CP�ROG���xe��`�'/sof�tpart/ge�nlink?cu�rrent=me�nupage,3�7,1 1  s�^��o��1631,�� ������l���4��C SDT_ISOLC  xi�� U��l�$J�23_DSP_ENB  H�|ai�?INC �H���V�A�@?�p=�̟�<#�
U��:�o� X������,�b�OB��Cr�R�����(�G_GRO�UP 1�H�>�< �^а�(�	t��?�n߳�� Q���� ��6�HZl��� �G�_IN_AUTO��T��i�POSRE�0�B�KANJI_�MASK��
KA�RELMON �xkf�Zry1J\@n����ӭ��	��(����� �CL_L� NUM�v��$KEYLO�GGING�P}`��h���LANGU�AGE xe�P �DEFA�ULT ^!faLGf��������9�U� �`��Zpy'�BZt� 
�Zq�Zp�#� ;���
�!(UT13:\��/ �/? ?'?>?K?]?o?�?�?�?�?�?Zr(9
O���; N_DISP ������������L�OCTOLc@ZqD�z~�Q��yAGBO_OK �o-d�4���1�1�@�R���O �O�O__,^?]{#��QY-V	�E�Ip��+�_O��B_BUF�F 2�H� 	�_���_�B(��_��� Collaborativ�V o%nmodovo�o�o�o �o�o�o�o3*<�i`r�SDCS ��ٟ��N\�_6�������'��tIOw 2��{ ��\���~��`�p����� ����ʏ܏�� ��$� 8�H�Z�l����������ȟ؟����;�ER/_ITME�d�i� {�������ïկ��� ��/�A�S�e�w����������ѿsG>�SE�V� 4M:�TYPE�X�9�K�]����RST/�uSCRN_FL 2�I�~Ч��������0�+�=�n�TP E��(�mMNGNAM�r��EP"$DUPS_�ACR�����DI�GI���U_L�OAD-�G %�j�%	DF_TB�IN���`�MAXUALRM"�mP���
0���_PD���  �COQ0�C/@��M��o�%�Aq��N�P 2��K �%	(������� =�O�2�s�^���z��� ��������'
K 6oRd���� ���#G*< }h������ �///U/@/y/d/ �/�/�/�/�/�/�/�/ -??Q?<?u?�?j?�? �?�?�?�?O�?)OO MO_OBO�OnO�O�O�O �O�O_�O%_7__[_�F__(�DBGDEF �{��q��T�_LDXDISA���i�9�MEMO_{AP��E ?j�
 �QhX	oo�-o?oQocouo�o0�F�RQ_CFG ��{��SA hW@i��chP<�td%�l��o�o�`��{��nT*?p/Ar **:JrhT= Ox�ohVu���� ��� �l_{�I� �`:�p�^�t���,(� Ǐ/����ُ���'� L�3�p�W�������ʟ���� ��$�&�IS�C 1�j�0p � r_l�nT�_��m_�����߯0�B�_MSTR� ����SCD 1��]�ׯQ�ӯ u�`������������ ޿��;�&�_�J�o� �πϹϤ�������� %��"�[�F��jߣ� ���߲�������!�� E�0�i�T��x���� ���������/��?� e�P���t��������� ������+O:s ^�������� 9$]�MKưa���ao$M�LTARM�b�:�g� ���P����PMETPU��PN���ND�SP_ADCOLx��P.CMNT/ %FN8 </'FSTLI]/N'
� ���.��a�/|�$%POSCF~'=G.PRPM;/�)�ST 1�� 4�b#�
L1XL5 \?j7H?j?l?~?�?�? �?�?�?�?,OO ObO DOVO�OzO�O�O�A!�SING_CHK�  `/$MOD�A�c�J���~YDEV 	�Z�	MC:wRHOSIZE�]N�UTASK %�Z�%$123456�789 �_�UWT�RIG 1�� l�U�oo���_8o����VYPvQ��T�SEM_INF �1�${`)�AT&FV0E0�=o�m)�aE0V�1&A3&B1&�D2&S0&C1�S0=�m)ATZ�o�dH4�a(o\�hAd�G���� �o��o�o �o�oe�������� r㏞��� �=�� �s�&�8�J���Ə�� �(��ПڏK��o� V�����X�ɯ|����� ��#�֟G�~�X�}�0� ��\�ſ׿�������� 1�����yϋ�>��� ��ώϘ�	���-�� Q�c�χ�:�L�^�p� �ߔ���N�;���_���p��|��rOD7ONERŠ/N����   ����P�SNIwTOR� G ?P[�   	EX�EC1TX�2^�3�^�4^�5^��P`�7*^�8^�9TY�� ��]���i���u���� ���������������������2��2��2���2��2��22�22*263���3��3i�QR_�GRP_SV 1�Ɖk (�A@H����T�=���>��}�{��=�Q��S�TR��ȉg!T�  �#��$>� �"]�)EW�fx�E�Q�\��,���ƓQ_DX�y^)#IO/N_DBP�]�!��� �@-Vn%X�w+�� -+X�N� (�!z-(+Y-ud1bU�/�/?Q�PG_JOG �����
(�2 � :�o�A=���?�(�I?[? m?61>�?�?��;�?`�;�0|2(��1@�O8O&O8F  �Q(��3STAT ��Z.1L_NAM�E !�U�@��!Defaul�t Person�ality (from FD)�"��@RMK_ENOgNLY�O�CR2�� 1��x����A; d�?_ _2_D_V_h_ z_�_�_�_�_�_�_�_ 
oo.o@oRodovo(� G1�o�o�o�o�o�op'9K �o r������� ��&�8�J�\�n��� ������ȏڏ���� "�4�F�X�j�|����� ��ğ֟�����0� B�T�f�x��������� ү�����,�>�P�b�t���(�<a���� ҿ�����,�>�P��b�tχkA�a@.���3?����(�P�� ���"�4�F�X�j�|� �ߠ߲���������� ����B�T�f�x��� ������������,� >�P��1�������� ������(:L ^p���?u��2� �  ����d �>�8F�?��0}�z�f  �����/�A�/#/�� (0m/4},�2�	`��/�/�/�!�1A�B�/? ?�?5 =@?9�**��0"�0C��3�  ��� (EW8C�  ä0��?��?��?O�?O:Oe	 >O%OzOeO�O�O�O�O�?�  �O�K�$�MRR_GRP '1�� QP(��"� � ��"P-P @D�#  @Q�E,Q?��A�@I�@U���O�  ;�	lXR	� �X � �P�R�Q ��, � �P�S� K�o���R��]K���K]�K	�.��Lv_�od�P@
�(baP0i�_�S��I�Xb�����T;gXb{Sў�]�3���b�1>�0�a�òN?v�?��=ڽ���?o0�o�bYQ�cT7�oUZ5�o } s��(p �  �  �8v�OV��U	'� � �trI� � � �L5�V:�����È=����u�R@��p�^2Q�BK2RD%��WyN� B�  'X�%aY`h�a`@e`h�mo#C�`���0C�`���m����"�_�_�XB� ���!��/=�q��Dz�O;��o_�pJ�o����R�����ഒА G4P��ŕ�zj1�K$  (�`?�ffW�����C � =�O��Q8�e�s�>L�p�`TQ�Z	(���P��ř�Q�U��R
���� x�Q;�e�m좢KZ;��=g;�4�<�<�ʏ�$��C��2S��<0?fff�?�p?&R��T@{=0d�?��p� ��"M�YT�O����ǿ 6��T'���� ��D� /�h�SόϞω��Ͻ��F� ���ϭ�"� ��C߽��v�ߚ߅� �ߩ���������<� '�`�K��o�{��� o_��=��a�*�u�N�0`�r���#��"�7&%�A��A���=���(��"���JH9��A���i�����q�� �����0�-�D1ſ0���� �l�`P�8,ȴA;��^@��T@��^5@$�?��V��P�z������=#�
���?��
=�G}�pm�{=����,��C'���Bp�����6���C98R����@\)���(��5pmG��p�Gsb�F��}�G��tE�VD�K.����I�� F��W�E��E���D��;.����I��`E��G�]zE�vmD���, �/P�/�/�/�/�/#? ?G?2?W?}?h?�?�? �?�?�?�?O�?
OCO .OgORO�OvO�O�O�O �O�O	_�O-__Q_<_ u_`_r_�_�_�_�_�_ �_oo'oMo8oqo\o �o�o�o�o�o�o�o �o7"[Fj� ������!�� E�0�B�{�f�����Ï@���ҏ����(��34�]�ء���P��8�N���3~�qml�~�`��5Q����`���ğ֟�������0���T�B�x�f���P�P������ӯ&�߯	�x��-������3� :�s�^�������Ϳ�� �ܿ� �9�$���0��cϙχ���Ϧ� ������� �6�$�Z�@H�~�lߎߴ߲�26���  B�R I ���CH"zm  @ Y�0�B�T�f�x���� H!����Т������l���?�� 

�����Կ������
 �e�w� ���������������+=O����������U�$M�R_CABLE �2Ք� ��T������� ���� ������� Nt6H~�� ���/��/J/ p/2/D/z/�/�/�/�/ �/�/�/�/?F?l?.?� �⛡��?�?��?�?O#O5O��*XO** �O�M ו	���������%%� 2345678'901�O�E �O�O��A���������
�G�n�ot sent �aJ�CW��T�ESTFECSALGR  eg���dZT3��A�lRà�����o��_��_�_�_ 9UD�1:\maint�enances.�xml�_
o  �B��DEFA�ULT��GRP� 2�yJ  ���A�ڐ�  �%!�1st clea�ning of cont. vP�ilation +56�Rڦc �a�o��+A@���o�o�*��%�ame�ch�`cal c�heck0  ��js�tq{�� �o�����?v�a?rollerRdv�k�l�~��������?qBasic� quarterCly�)�;��j,[��(�:�L�^�p�7yMXI����"8������ǟ�������*�<���C�f������㟸�ʯܯ� ��?qOverha�u�����>� x��H�O�����|�������Ŀ��$m��O ۿ��k�@�R�d�vψ� ׿���������� *�<�Nߝ�r������� ���������Q߹�8� ��'�߀������ �����M�"�q�F�X� j�|���������� 7�0BT��x ���������� i>��t�� ����//Se :/�^/p/�/�/�/� �//+/ ?O/$?6?H? Z?l?�/�?�/�/?�? �?�?O O2O�?VO�? �?�?�O�O�O�O�O5O �O_kO_�Od_v_�_ �_�_�O�_�_1_oU_ *o<oNo`oro�_�o�_ �_�oo�o&8 �o\�o�o��o�� ���M"�q�X� �|�������ď�� 7�I��m�B�T�f�x� ��ُ������3�� �,�>�P���t�ß՟ 矝�ί����e� :��������������� ʿ��� �O��s�H� Z�l�~ϐ�߿����� ��9�� �2�D�Vߥ� z����ϰ��������� 
��k�@�ߡ�v��߀��������W��	� X���-�?���B `�n����������� ������"4FX j|������ �0BTfx �������/�n� Ў�?� ; @�� L�G/ Y/k/��3/�/�/�/���*�/** F�@ h�j� /?�&?8?�/\?n?�?�?����]��/�?�?�? 
O�?.O@OROdO�?�? "O�O�O�OO�O__ *_pO�O�O6_�_�_�_ j_�_�_�_oH_Z_�_ Jo\ono�oBo�o�o�o�o�on����$M�R_HIST 2��f�"p� 
 �\6�$ 2345?6789012:t�o�"19/�� Z�-������ E�W�i� �2�����Ï z�珞���ԏA��� e�w�.���R���џ�� �����+��O��s����<�����pSKCFMAP  f�%p�"	q������ONREL  ��"pڡp�âEXCFENB��
أ��%�FNC�,��JOGOVL�IM�d"su�âK�EY�x���_�PAN�����âR�UNh�x�âSFSPDTYPL�<�£SIGN���T1MOTj���â_CE_GRP7 1�f�ڣ*r ��/vσ�cϠ�Ċ� �ς���߸�%���5� [���6�xߵ�l��� �������3�E�,�i�  �s�����z���������áQZ_E�DIT	�ԧ��TC�OM_CFG 1��Э/�|����� }
]�SI �M�B��������� �������W~6�T_ARC_)���W�T_MN_oMODE	��T��_SPLz:�UA�P_CPL�;�N�OCHECK ?�Ы ��  "4FXj|� ������//���NO_WAIT�_L�R�=�NUM_RSPACEͯ�H�/�'�$OD�RDSP��7�O�FFSET_CAqRH���&DIS�/��#S_A� ARK�	�S�OPEN_FILE� ���S����OPTION_I�O����T0M_PR�G %*%$*؍?�>03WO0�M���p�5�i ����0��1�	 ����3�f����� RG_DSBOL  wڡ�@/ORIENTT5O���C��١�A �"U� IM_ED\7ע�� V� ?LCT �+�d�t���I��d�i�C_�PEX� �/�DRA-T� d7��D� �UP �N'p��`�\_n_T_�_�Y�o$PALe��M���P_POS_C�H0_�QRAM2�F���x;���C�@I %o7oIo[omoo�o�o �o�o�o�o�o!3@EWi{���2o ������(�:�L�^��������� ��Џ����*�<� N�`�r���������̟ ޟ���&�8�J�\� n���������ȯگ� ���"�4�F�X�j�|� ������Ŀֿ���� �0�B�T�f�xϊϜ��p<w���������� �0�B�T�f�xߊ���kA�a�r�#�� �y�P���ߞrP��� &�8�J�\�n���� �����������"��� �X�j�|��������� ������0BT f5�G������ �,>Pbt�������r	F�!���KBd� �/,-/N/\'��@F#�/��/�/|!�0��'�/�/�/�/?2A�'?9?�(��0�?�<�r�%	`�/�?�?<�?�1:�o�AO�O,O>OG A� � UI�(@!@!�p"��pY$��C_�  ���P�PoFC�  � �@�/�O�/�O�O___P_{%	T_;_�_�{_�_�_�_�_?� � �_k�$PAR�AM_GROUP� 1�#0(�#K�� �2� ۷ �2Fa @D�  ZaeFa1?�pa�qC4\cZa����_  ;�	l�rb	 �X?  �`�b��a �, ǀ ��`�c~0H�����b���H����Hw�zH��\�o�",t~0B�  BqzaJy<Ys�3��rr�A>�@sq��ew	�0�B\�
�Ѵ9��1K�^G" ��rsa�jG�epE�� }:��B����0�  �  ��R��_p�u	'�� � ��I�� �  �<bEv=��Ͳ�ċr@ڏ��~La���;Lb^�?�wN<@\�  'r�~0C�p���@C�p���0���������B�o�oxB@
�A�EM�2��1Dz�_U���y�d�����r��Ƣ��΢А� 4PΒߥ�5zȀA?"����p?�ffm/�"���C �0W�i�q8�0���>LԀ�naz	(�0��Pĸߩ�a�e��b$���� x}1;�e�m¢KZ;��=g;�4�<�<��/�>�c��Lc��R@?fff�?�?&l�t@{=0~�?��� �9Bg�sd�_������ PǦdA���:�%�^� I߂�mߦ߸ߣ����� �����6������/� ��+����������� ��2��V�A�z�e��� �����+��o��W� {�D��hz��=�c�<�M6?�A���[�W<'"��d^I�;C6�p2-�%�3?��	p��/� �x`1�@M$D1��J�������!@I��R,ȴA;��^@��T@�^�5@$�?�V�+~0�z�ý��=#�
�� �?��
=�G��F-�{=����,��C'��B�p��� ��6���C98R����@\)��(���5F-G��p�Gsb�F��}�G��tE��VD�K6>����I�� F��W�E��E����D��;6>����I��`E��G�]zE�?vmD���F/�? j/�?�?�?OO=O(O aOLOqO�O�O�O�O�O �O_�O'__$_]_H_ �_l_�_�_�_�_�_�_ �_#ooGo2okoVo�o zo�o�o�o�o�o�o 1AgR�v� ������-�� Q�<�u�`�������Ϗ ���ޏ��;�&�_� J�\���������ݟȟ����7�� (�!3g4�]9����j��"�R�h��%3~�m8����z��5Q��į�z���ޯ��!���
�
�J�8�n�P\�����P*�Pľ�����@���#��<G�2�����M�T� ��xϝ��Ϯ������ ��/��S�>������}߳ߡ�������� ���,��P�>�t�b� ������� 2P���  B�lc�C%H< zl� @s8��J�\�n�����������������#?M�, 
$��#��%� � ����
 ��� ����!3E�Wi�*���������U�$PAR�AM_MENU �?
���  DE�FPULSE@��	WAITTMO{UT�RCV�� SHELL�_WRK.$CU�R_STYL��,OPT"�"/P�TB7/1"C/R_DECSN���@� �/�/�/�/�/�/�/? ?$?6?_?Z?l?~?�?��SSREL_IOD  �ޱ��5�USE_PROG %�%�?O�3CCR��2ޱ�G�_HOST !Ʊ! D]OJM_�DA5 �
��Xe. ��G���=���7���C�vETհ'O�C@ORA��C�OK_TIM�E��60E�GD�EBUG�0��3G�INP_FLMS�K_GYTRV_GWP+GAtP 7\���[�CHU_FXTYPE
����?�?o5o 0oBoTo}oxo�o�o�o �o�o�o,U Pbt����� ���-�(�:�L�u��p�������IUWOR�D ?	�
 �	RSuPZ�P�NSX�$��JO�N![�TE�@��COLXŹ�D��WLV�0 ��C��0E�d,QTRACEC�TL 1�G�� ° ݰ�ݱ����DT Q��
�ِ��D �� 	/�� �M �Y �U ���������I K&�1ܱ�1��N���10�f�	�&�ݰ����6�����ʯ ܯ� ��$�6�H�Z� l�%�q�������ѿ� ���	��=�O�a�s� �ϗϩϻ�5����� %�7�I�[���o�aѭ� ��9����ݵ���a�� ���0�j�|���� ��~�H�Z�����0�B� T�f�x���������� �����.�*<N` r������� &8J\n� �������/ "/4/F/X/j/|/�/�/ �/�/�/�/�/??0? B?T?f?x?�?�?�?�? �?�?�?OO,O>OPO bOtO�O�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o o$o6oHoRe&to�o �o�o�o�o�o�o (:L^p��� ���� ��$�6� H�Z�l�~�������Ə ؏���� �2�D�V� h�z�������ԟ� ��
��.�@�R�d�v� ��������Я���� �*�<�N�`�r����� ����̿޿���&� 8�J�\�nπϒ�ho�� ���������"�4�F� X�j�|ߎߠ߲����� ������0�B�T�f� x������������ ��,�>�P�b�t��� ������������ (:L^p��� ���� $6 HZl~���� ���/ /2/D/V/ h/z/�/�/�/�/�/�!��$PGTRACELEN  �!�  ���� ��&_UP �����!1�)01"0�!_C�FG �!5T3�!
"0�N4N4�h?s70s:  ��s962DEFSP/D �A<�!0��� H_CON?FIG �!5	3W � � d�4M�2 �!�1P�4؅1A� �� IN~90TRL �A=�a18�5 APE�5��7�!1N4�1��9LID:3�A=	~|ILLB 1��9_ �EB�0sB4�Cs6 H��G�OEu? <<7 �!?�[-_ _%_G_u_[_}_�_�_ �_�_�_�_�_)oo1o_o|j�B�o�o�o�o�_�o�o�o5{IG�RP 1��L��� @A!���4�I��!A �C�u�C�OCWjVF;|S0��4`�1�y�y�1�0��@04_�A�~´���{B�/����E��/�i�{�&�B3�4�����Ҏ��#Pj��׏�ӏ�F�1� j�U��y���u��ӟ  Dz��R1 ��>��N�t�_����� �����˯���:��%�^�I�����)���
V7.10be�ta1N4�0@��*�@�) @ߺ+A �2?���
?fff>������B33�A�yp0ͳB(���A���AK��@kqxq 0˱˴̱@�+�=�O�a�xqp�����1l�ϥϱȿ���R�fh����oB�!x�Z�t�z� �����%��p߻��4	/rqBu�N�!5�� � ����iA����wӛ B�0B�����B)H%��� �r�&G��Y1�W��x[�x�߁��߉����`0z�hB���1������A�����A�ff+�ia�D�KNOW_M  �~5I6�DSV ��:BS,��� ����D���=�!��} A��*SY�STEM*� V9.40341 {�1/17/202?4 Ac� h����@MSq_T �  � $MAX_PYLD�0�$AXISIN�ERTIA   	$PS_��7�L� � �M�OMENT��_Ơ SC� � �WT�	INR	 7 MN.�CL(PLD_M�ODEDUMMWY11�0b2j�� MR� � {$�_ENB0�$W}��A�NGL]�@}A�A0�B��CCv�DD�ST_��,
$COMP_�SW�0�XY_LO��Z%� ��� �� ��}�AYLOA�V7#_X=*Y=*Z=*UIJ+IX+If#I�0�DISP0��4� _RES_G�� | 5*S�AV�� �)5�+6��%��&��&��#EL�� UL0 �*V�!  �@�$A��PMON_Q�UE�!A@$Q�COU/!�QTH&� HO�r0Hj� [IS~3UE]0U�!O�PO�@�!�7$P[BU���OVERRUN_�TO�� ODA�TA�!
@�6C���CUR$DE�X�PROGRA�#� � 2NE_sNOD�5ITPCޟ0INFO�! ��0�;/A��31O�I2B	 (0SL?EQ_NUMFC2@�YP]qB�6�1S_�EDIT�!
 �̊ K_�@kC$_HIDE_� U�G��HAUTO� �EC�OPY�A�0�Lu�$RMV_MAN��@�Kv@�3PRUTؑt��NF�0UC�H�G�21T�"RGwADJ�! h� kX_� I�1$  �]V ]VW[XP[XR~[XSPEED_MP��NEXT_CYuC�GSNS_�3�� $ALG�O_�0�NYQ_oFREQ�WI�0�wE�QSIZyC�1L�AS�Q[Q#�PkEC�REATE}3�0I�FY�6NAM]�%,d_GSSTA�TU� S�7MAI�LTIJ`p1waEV<."�LASTwa�!��TELEM�Q =��ENAB�`EASI�ap1��� �bkA��f�RO&0ATI@$�R��u1� rAB�1<l`�0D_LV�a$v�BAS~a$v�`?sU�PD_�0~`$�<qXwRMS_TR`s�� ts�SP}3`�aXt�B�R#� �	�b 2  b�	��wbr�w�rZ �br�w6%�RARN_DOU�3��IN��TPRE�-P aBGRIyDA�3BARSjF8P�c�bOTO� �!W �1_Hd!�P�o�/�O��T �s �POR�3������SRVL`)�����DIRECTA_iҀ�u�3�U4�5�6�7��8Ё�1FXq�1~�0$VALU?s�GRO�2�d� *AF>�U� !�e���1��Na�0i�RAN��v�^aR�@wAp1?TOTAL_{d
p�ԒPW�SI7��R�EGEN���3X�ex�3wE91��X0TRKsib�_S�0K�����cV[Qii�ukaGRE~c;�w1o2�2�@n��V_HX�DAX#k���S_Y�Q��V�SdARX 2 })RIG_SEn3�U����e_�0��C_�c�$CMP��D�EV1 ݠ#�I�P�Z�DF�HA[NC^1� 
�gq^byC��INTπ�QGF�3!MAS�KZcVpOVR}3P�O0;�t Ma�L�OV�Cbij  M�:�� 4f0H�jF%�c��OPSLG��Q�r@� �V� Zѐ|`S��d'�U��7I�P}�V���`�T$1O����CH���R!�l �r4 *$�uA��J ��ACcIL_�Md��Vr�`�T!QX0�3A_pC'6�5V�C�P_��~`�$�M;�V1:�V1�H�2W�2H�3W�3
H�4W�4H��1i�r`�1u����rIN��GVIBh��2�U2�2�3�3�4�4� #Ԫ"� �0������������;PLc`TOR\0�p��Գ��BRK��S�3�� ����� �^2d� MC_9F{0� 	e@��(��g�ǐM+0Ig��� � E"'�� K�EEP_HNADED	�!K�)pU�C*!�L`k�o�
�� l�O Q1J��@��l�l�l�REM��k�{a���������UHdek�HPWD  K��SBM����COLLABZ��2�ő2b�J@IT�P��N=O9!FCAL�ē�DON�R���$� ,0FL�~aO$SYN�yM�����Q�UP_DL�Y�!sDELAh� |a[bY� ADX!�$TABTP_�R��QSKI�P Ĩ��0O0�u��r� P_�0�2  �0�� i%u %�$�$�$,��$9�$F�$9!q�{RA�3 Xܠ�i���MB��NFL#IC�3��PU���7NO_H� ���A^��SWIT2R��_PA @G�q� �!1b�UdpWJ�O�:#ߣg�NGRLT� �1{Q�K�M��<!�pT_Ja&�r�AP�WEIGH��3J4CH�0a$O1Ru�a$��OO���bD�a_&J���q�SA�!��#�(OB�`�Y$�)p!q�qJ2�_1�EXJpT�S71#A p171JPG�71AG����RDC��m ��@R����R!a��q<���tRGEAD��`���FLG���0�(�3�ER��rSPC�"C�QUM_70��2�TH2N2@�17  EDo��R   D `�\�)-p2_P�EC�S[��q�PL10_�CbGPE�� !UP$K@мp�3 �v����A�4�P�1���uKA���CE`���r�-s{�Fz�&@" P>,@DESIGbB�uVL1JI1WF�C	W;10��_DS���|��;�POS11w�# l<�r�N�x�1#�/AT��"��U
8�RIND����}Q�SP��}Q`"�rHOM�E�R NU2WR$ ]_o_�_�_�_�_`PS3WR%�_�_�_o"o�4o �OT4WR&�Woio{o�o�o�oFg5WR'�o�o�o
.��OT6WR(QcuP���Fg7WR)� ����(� oB�Q8WR*K�]�o�����䥏�US XQ+  ��PS��0C��<K ��, T,@]�Lʖ]�IO��}�I�:��OK _OP����x��1nCPOWE�я- G�x U1#�P@�YP.sؒ�$DSB3�GNA��B� C@��BM=Ic�/ ����)�1�0�7 $T�P ɣ�෰WAI4�@>g KE� �3�Y1�X��H�S���)ޡNEC-� � J��2�AL1ƦAƢz�1t�OT�S�1DLV�IC����W@;QI߄SBN�%h0n�PEA?�0�p0���>20�ACC�� ����H��5H����g1 `�]�UF" �[�UTOOL\�M�9UO�W2NC Rq_��s�AND÷��b���2w2BU�FV���M� R_V3RS���IN�2@ ӰH�0����(�_2 <�>���4�,�|3Ǿ�A 30<��q�|�1 h0S2;32c�3 �y0ͅ9x�D�ICE< �cPE@�  IT���OPB7 �FLOW�TRa ������CU��_�� U�XT��4 TER�FAC�İ�U����rSCH��4� t<��B����!�$FREEFRO�MW���GEX I�	�UPD"�iB�1PT>�p%EX��g�!�FA%�C�8 ���P�6�5 &
̈; A| �ى�0�EX�IO#рRYY����_O��P�ь���WR���Dp�1/�D��FRI,�z@7 ����j⢶j��MYH�i�+�GT_H_VTEY�I�A���P$CPӰ��UFINV_SP��H��RGI��f!ITI� ��X�����G2��G1���@��� ��PRE_���<!DI7"���#��t����ʐC> ��9�u�ALAR�0q$��Z�J�� �T�ҭ�$�� o@% $�6�6 @n��0��P�d��"��$�A �� B���7X �;"M��CT��H@�@�0���Դ�G�3AW�m��= �D� ��Kq�� ϡ��xA���� 26ʀH)�WP/�1;�*�2-�2�3-�3;��	- <��	I������!�$VϠ��V��V3�����U�7�8w0 #ֿ=�V2c��¹�e�4�S�1E�0c��A����A����@�PRQ0�pS�1�!qܒ��f�9 
P��1+� 740�� 8 ʀ��:��@FR
�@�ҽSʑ: ؠR��!1�Bo�U��°X���S�ұL��NB�"T�H�ԐI���@F�ER��4C�"IF_���&I-��#�� GA1(4�$9ĵ<67_JFE7PR�AIP��RVw; g $�A��  �BVALU�1�0j6zC�<Вx� 2; ��SCʒ=
  �$G�4A�2���4qT�@�#�3DSP�6�JOGLL���Y�P`0�5��!�3^@AXt�z�K}�_MIRAd!D9�MDBEAPc� E��&�1SYS�8A���1PGwFBRYKU��NC�0I�  �B.�B�2��qD{��3;@BSOR���3s�N�EDUMMY166i�נ����z�FC�_OVRi �� �LDRCOIRW�NF�VF�!lV�0OVESFTZ� WSFpV��%C=���X����CHDLY�G=�OVT���0Wb��M���U@RO����A@_� �  @�d���VE_���OFeS��C�0Z�WD8Q��T4Q�Aق[E�@TRr��_�9�FDO[F�MB_CM��F`B�0BL�?�hb�+$�V$�o���3PRGig|HAMzC\`AЪe�R�o_M�`�9�x��PT$CA�09���>�T$HBKs��&qIO-�u��O�PPAz?q$yOt7u��e���RDVC_DB��q�!���p�R��"�u1�z�c�u3�v�PATIOF�0�QqU2��0x�CABY� ,�B�= �S��h�0�_
��&SUBCP	U��Z�S����Rc�d�t��S�p�dՒe1$HW_C���䅇�A#� �$U�NIT�D����A�TTRI� ��Z�C'YCLC��A�rLC�FLTR_2_F�I4
��s��LP�K�4�SCT��F�_��F_��8���FqS���b��CHAF�� �y��b��x�RSD����������7p_T��hPRO�p@c��E#MP��@�CTf�wa��g����DI�О�$RAILP�/�MF�0LO�@���D7i�`��v��u�cPR�p%Sw�T�X�Ctq��=	�SFUNCd2��RIN��s��AG�w���RA��t�R�Tp��D@	t��WAR53F�`BLq�ѤAʫƁͨƨDA갡��ѣʥLDd�P��4�d�!Q��3�TI��S��1� $/ RIYAHѽ�AFD�Pm�~��P��� �����MOIG�CfDF_�+��Sp���LM�cF�A��HRDY�ORG8�H��wQ'��>ҵMULSE+��#TS����JZJ6R�KWF[FAN_AL�MLV��R�WRNY�HARD�@s�����J�!�2Q����1�E)_�P��U��Rk��?TO_SBRvr����0�ʥ�vs���MPINF� ����)�n��REG.�NVq���ӚFDA��RdFL��d2$M��%R�d�`� `�g�CM� uN� Y��NONI`��N�DEVY�j�s���� �I``�1>� �Y�$���$Z�� �2�1�0?o, �oCEG���3P�ѝ��t�E29pi����|EAXE�7wROB�:RED�6�W��A_]��CSYЯ@8�p�S��WRqI�P慀STR�5(���@*PE���0�C!3O �@����B���Qp��]��@�`OTO�9�0�PARY�3�0!��t�1AFI�@,C?$LINK���!J'�c_���Q��:�N�XYZw�Y��2!j�OFF�P&��N�B��B�0l�`���q̐p���FI)Р��w!R�Dl��4_JA�2(R3�;q����4��9!�TB���25C��kFDU��E�354�TURT�XZ�n���X��pFLm�P��� p�x���Ca 1>�0K�pM�$\3�S��S�%cORQɖ�1����84��@10ð�<p�#�1#�QOVEX�"M,�01��r��r ��q��o�p��o B5q�,����!Y9@� �r01jYv����L��1ERA �	8�!E�Pn0D�9$A�� ����Ē����AX�S�2�����(� �%���)��). �*e  �*�@�*3��*3�*!��*1���&���)���) ���)���)���)���) ���)��9��981,9x���~%DEBU}�$x�����1bJ�CAB�q8QRVp|� 
B�s!/E ��;G��;G.;Ge;G �A;G3�;G3;G!ኴp: �����LAB��qy��sGRO��4}��`B_ґ & ��͓�����FQU�� VAND� 8�.$ �qS�1!��]W �a�����qX��X�R�NT8d��S�PVELؑ���Q��X��͒��N�A�a��h�C��0%TRQL��Vvd����SERV9E�P��@ $��n�Q!1`POJ�}�_ĐT9�!� b����A  #$Ub `�
Tch�2^`Bbg��2Aseb�~�_ C lT ���ERR���Ipp�P��aTOQ���L<��$���fĐG�3e%<�|" ��VaR}E� D ,/a�we�`B�RAq �2C d8rfs�uj` E��$�fג���"
�TcO�C��`F  >�kCOUNT��sFZN_CFG]aGG 4��%���T|# z��q�3�Q�ab`�Ѩq^��H �,@Mz��+�!���oz��F!Aq����XX�5� ��a"G�4d̀X�9Pz���HELAЭr�I 5��B�_BAS|#RSR$�`�R�S<�L����1w��2Ċ3Ċ4�Ċ5Ċ6Ċ7Ċ8w��RO�Pq-�Q�3NL��@AB@c
�n��ACKFINfpT_U�U��	���T��_PUX~�e�OUBcPà%؁�v�����y&TPFWD_KcAR�a-Ѻ`RE?d��P#����QUE�$�f YI �~���I U�C��O𲓲P�O�SEM��G�EAȰAn�STYc�SO2�DDIo����C�x'_TM9�MANsRQ��O�ENDD�$KEYSWI�TCH��Ǒ���H}EI BEATM��PE(�LE�bґ PJ��UƓF6�ǒS���DO_HOM��Olz�W�EF9PR��P�rj��U�C�O��<�`qOV_M��E��OCM;�EAo�P��HK��GJ DL�&��pU�b��M�ᔒ<FO�RC*�WAR�1�D��OM� K� @�4���U��P�'�1�g��3�4�QQbkpOא`��L<$r%�UNLO���dmb�ED��  `��@HDDN]aM �d`BLOB  � ��E�uN <�NЉ�y"��MSU�PGB��CALC__PLAN��1���AY��{�3��tO '� ��9 PI`$ MѠ��5�B����Q-�Ml��C���ƹ�d��SC�eM�ЭQ�` �aѹaQpt�Y|�Z�|�EU�,��[�T�aU��bе�PrNPXw_AS�rP 0���ADD�p�q$S{IZ|!$VAP~uMULTIPD�����A��Q � $����F��𐲁�М���C�`G�F'RIF��fpS��	��J�7�NF��ODB�U� �PH���?fCM��$@�1�C�t���.�q��)`R �3 ���bTE�,.3SGL�T5� �&�p��C��ST�MT�5�PSEG�@�5�BWY�SHsOW=���BAN �TP����A�,0��7A$�=�_CT�>� S e t	p���`��A�LI%b��OPEN�F�Q�q�WA��NEW_L�Õ���B�����q��RIL;N_�BLK�P,1P�- -EXp-;SY�IPE��q�Jp�TCz�B	�P�t�Ʋ�� _BUF�RNW�� PrV�+ _G�rT 3$�PC�@gp+#�!FBZ��P�SP�An�����VD� �rU�� ��aA00 bT#�+'�+1�+T;�+5)6)7)8)9)A)��+ �+�A,��+� ++0�51B���\U1i1v1�1�U1�1�1�1�U1�1�1�2(U252B2O2\U2i2v2�2�2��`�(�Bp�(�U2�2�3(35U3B3O3\3iU3v3�3�3�U3�3�3�3�U3�3�4(45U4B4O4\4�9U4�94�94 I4IU4�4�4�4�U4�4�5(55U5B5O5\5�9U5�95�95 I5IU5�5�5�5�U5�5�6(65U6B6O6\6�9U6�96�96 I6IU6�6�6�6�YU6�6�7(75U7B7O7\7�9U7�97�97 I7IU7�7�7�7�Y�7�i7��VD�_�UPDV���� 
��V��W x $TOR �����]�O�p'�t��t?Q_CURR��ZԣAXO�ҰZ�S�}C"��'�_� 1����YSLO��X � �Չ▣r���,��p%�^�1�VALU h�y�̖�q��FO�y YL����HI��I�?$FILE_-��ƽ�$G��M�SA�VY h�p�E_BLCK��#�-�>,�D_CPU<���@<��к�����Y���k�R Z �� P: TO(�6��LA|SR���\����RUN�Gŕ ��ɑ��ʠ̕ꑷ��¬�Hด��� ���T2e� ��[?  $JP����^�TPP_EDI|���T2SPD,��\4�X�S5��� ��DCS��G�q�] � $JP�CQ�'�
7�S��C���C��$MDLf��$}�éTC4�&ŧUF�pĨSF�ĨgCOB����T1��QT����^ ���Q��5�����?TABUI_����y_�� ]��.��^$��A���LB_AVAIYР� �I�`�p�$SE�  1�DGE_ɐN��¬pA* !N�Ň�Q�E� ��$����_}�.�_��1�wELE� ���SCRN a )D��òB�T!ò4�r��pNOd�V��@�PRIO�t����Ӳ_MP��b \@�pf�b ����M��JD G� U���6_�SPS7��NѰ|�z
�E̲�TBCD����c ̡C_B�RK2_MG���H�!�2dW��e�B����,�FTMh��rf�2 �DC���C�б�`��x�THD}�u��ԩų�R�{$��ERVEk����x����� BC_�$� 2c 	3� �_AC�� e�X -$�LE�Nk��x���RA[TI-�$N�W���F1�ׄ2U�MO�4���@��ERTI�A��}��t���D�E��8�LACEM��wCCp�#�V��Xp�������TCV����TRQ�#��@���G����J����p�� J��������29�;�������JK��VK�k���x�������J0l����JJ��JJ��AAL�� �� ��e4 5��$�N1*� 6 �����t�α�v��CF��f `�pGROU��v�f���N[�C�� REQ�UIR��$DEB�U����L���e���б �SGI�gz��e�APPR��YC�#�
$=�N'CLOr�S��)���
 �ARA[�h �"�2���#��d9�1�GR�xL���xy5�wNOLDw��RTMO+���hJ�@�P���� �����#��,������7�8=�nI�i�� ��5���xT'x�b#PATH^'�w!m#w!:�s#T�h%�NTe�Aj��6mIN�UC��b�Z� CL�UM�(YW���p�!Á���*���*��� PAYLO�A�J2L�pR_	A�75L��C9?139�O1xR_F2LS3HR��|1LOD4�!p}7�#�7�#ACRѠ �(�0�'+4��H����$H:��2FLE�XC�$�j Tr�MR4���kDh(4�Π:KP� B7�Ѳ;BJH�k l�W��i�������_FUNr��W�E��j 	jA>�l :�,� ���GT/�ѱ�8�J�\�F1QaUuWk�}� ������RE���� ����)�;�M�_�|h �da�����c��h����H��Q��T��zaX�� ��X���W��Ju#h�� ���� ��#,�>Pb	��BJum � ����Q 	ĐT��k�U�0���a���J�yAJE�C3TRҊPTN)�\���HAND_VB� BjAOPoEn M$�`F2x����M��BnRo� $AdR���0� H� FA_.2h)DU�qA�A�9Bz��H@�D�IB?I̲XAGR�XASTЖXB�XAN�DY �0xD�k�A0�s7 Qs7�127���d;Pp�P�%%% %)%p2%;#��oEp ��D\" �Q��6�OASYM�%=p�B£$o�P�-�1�/_SHi�'�$�P�Ԉ�/??%?73J><�P:p��o9�T_VI���,�6=�V_UN!I��Q�ss{1J��j� ��j<nĥ5{ğƮ=�k��9��?�?��+sh�4 C�E�CH�?qP |A���fTO/`PPp�VP��B���aR!PP�@�`eF�i�e�I�_�5�!P�І�EѮ �RPR�OG_NA�Q$>a
$LAST��c�CAN?P3�E�XYZ_SPA�U���)���}@��S"м���E��@��CURd�FI�R����IO_TY9P�cJ�IND�G�.�X��E�p � H7R_T�r͂��"��P��cO��B���s �pr�J� � j�� ��Pz���P�l�p �P�� t �� �ME�QМ ����|�T��PTDҰ]���p�t|@���"�=�1�TӰg~+�DUMMY1{q�$PS_�PRF�NPg@$x���F�LAw N��%�$GLB_T������3�p LIF��uc�R �s�OW��\�d��VOLw�.�&��_2�!g�2;!g����b����+�TC~yQ$BAUDBQ���STBV�s�A�RITY<D_W-AUAI!	C��Q�OU�1f�	TL�ANS��`SZ<(�BUF_��@p2`�J�CHK�@�OCESUQr�JO�E���� ��UBYT�B�A �"^$:m$����CYܸB��SCR�� v .�E�P�P�RމPLUG�����-���w L �$PWUP.�k�P�Wt��L�Xk�EE�a�fIU����g)���PR�����x 8�0PISN5d�%6*7d��o�����yL ������CHX��pu(OPEPNS@���e����'��
e�2#�#-e�9 e�Ae�O�"]�'3s�#�	�M1�	\7 �M1�M1o��q����P����z XX���pASTw����SBR��M21_�KХ`T$SV_E1R���5�3CL���2eA�POj�|�GL4��EW��{ 4 m$]�$a$�$W0C���ჯЩRy�FUE|��$��$GI��}$A @CI@J��}�jG��};�z��EsFNEAR�PN��$F�I�PT�Ѿ��P�J��R�X� ~�$JOINT-q`��A�MSET��  "hGE�E�Q*�S1��E|+�����  �P�U�Q?���LOC�K_FOL���B�GLV��GLdXT�E��XM��#QEM� w��R��OP$cUS��@-p2|���IC�Q}yR�TP�Q{��1CE�p|C�P $�KAR@aM��TP�DRA@�T�AVEgCLEj��DIU�Q�~�QHEVPTOO�L��+�#bVI,cR�E`IS3q?e6L�qn�CH	P9�*�CON#�<%#8`I0�� @$RAIL_�BOXE-qG $R�OB�ЁR?��1HOWWAR���au�jaROLM���e�q�gd�b � :�ǀO_�F!�!��HTML5e�3�Q�܀.S���@\a����NAC��e�TP����BSLO��A�`�A� ��� 	t���U{|�f�u�OPVrPOXq��I���TN� 8b�b\a�ЮQ|/p��ORDEDTP�9�Np�@XT�pQ)����M� ��� D ��OB��j�TP��w�q�S���a |�YS�qADRk�|��|!�*� � ,πN��$A[Q��Y����C_|�VWVA>�� � ��B��"RT��$E�DI�ѡ�VSHW�R�`�1�4�0�LA�aH�Z�NBՃSH�EAD�����Ǳf��KEa[�CP��.�JMP	�L���oRACE����p�N�I�PS(�CH�ANNE+`)��7T�ICK,c_�M���/�HN�1� �@�pL��CP_GqP�f��STY1��haLO�����(-������pp
�Ь�S%$~���=�0S~�!$`�� �N�M�9PB��SQU�Pޣ�LOO�+�TERC�!���TS4��C r@��c�Dp�r��a�#��IZ����L�t�����4щ P�ʥ_DO���X�X� S��AXI��b�Q.�&�T�Њ��_�FRE3Q_`)�ET*���$��\ AW��0
�`H���AT�J��h�9�� �BSsR_�1F��lj���p�RQ�C����0���B�ѳ�V�ѥ�NOLDӹA]�A��tO���A��AV_�Š�ʿ��D�D�(�� <�J��C�C��)�C:���CYCn`w@��n`_"�������o�	z�SSC��� � h�`D1S����u`SPq��AT'���ˡ��X��d�ADDR�$�T =IF�ӥP_2�CHL2!�I�0L1��TU�0I�� ���BCUO K�ApTV
9RI��J�dX+�M�*�
�Z
�VgqڡNF�� \��x������@��C[Ë�N�p�ڀv�2���TX{�EE�r���+ }PICNACy@I�Dv�8+�+�
Б T>��0 ����0�0����{#���䥀RR�A(���|����  �UE4�G� ������S	AN)�RSM���U�p�T�� �THRS_ CC ����#�>���+��CIR��}� 2�vD�UE��� ����b�� GMTN_FLg���0�q�A^tBBL_l`W� NF�� ����O=A��LE[���`�����RIGH�RD<�4Q�CKGR� �T�pWIDT�H�3��"%FLA�G���UI�`E9YpE�� d!@p��`̒� �aBAC�Kʑ�b{�1u F�O�q�LABձ?�(u I*PMR$U�R�a� �@T MEN�H�� �"� T!_�L2�؀R�OR �3rh3� P�Ob�F�%���GO0U��,9R]R�aLUM,�&�K�ERV�q��T P|�@[� � _��GE��AI��r�LIP~G�EQ��)�@������V`�5�6�7�8�O�������@
�te1�2GQSv�@�SUSRDO� <��� UoB̞�oBFO��oBPR�Ig�mv`��} TR�IP�am�UN,� 4��f@�� 略a���R(��0� ��H ��G ���T�`��M1�"O	Soa�&R.����#(a�A�O1C8N2��7%0�#U�A�?+?p9����#OFF~P*
О�A3O�0�Pќ�`�4�4��`GU#�P�1Y��3���7h�SUB�� �E/_EXE3�VG��#�WO�� �`0��'�WA��H Az� G�V_DB*CHB@��H T0�������A�`��ORl`rERAU��sDT�IA�XAy_��4�� |���A�OWN�P`�$GSRC��H��D~P<�E��MPFIÔw�*�ESPơ��a�:e [}aWHb��C����G� `b0B`���n/�COP�$�� _�@r�lQhqsU4BCT
A&SAHb� �~��b�� ���SHADOW�:c�Q?_UNSCAc�S�@�SDGDaa�E�GACfS���V�CͰCY3�� ��b"��$`EAR��/l-�t��Co^/eDRIV��5�C_V��Rd��a�D)$?MY_UBY($7d��3���.�a�ہ�h4Q�bP_�PÔ�bmLЫBM��$W�7DEYF�EX�p��wUMU#�X��"t�cUS���x _R_�l2m 
���m1G\�P�ACINg��RG �A[tqrw3qr63qrH�lQRE�_�1Y�8cqr
Х ��^PeGw`P,�p d	R 0
Цc %��I��2	kR�RE.sSMWip_Ajq��#s��O>!Q�Ac�*���EE��Uې� Z�� VcHK���"B�`B���'���s�EAy��}�@o@*�0bMR�CV7�� �wO*�Mo@C-�	���3�s��REF��܆Æ ���hX��M ���@Њ��4�Æi�_�@�j����S w�c�z��AM1b}�� �@����r��Y!�el��OU�3��r1�7c g��u��2���0J�๠���*�������K�ULW��f+PCO��fP�p�NT&SS�4RR�^�5!^��L�c���c�����5!�VG�R����� �$����O� ���BVLO��$X�������I�SY����QDOx`EQ&#��c�2�PIX�w31�SZ#��d^��d2�H��`ВS1�Q��B��SI b�l2��������}�f� � ^r~�a�Ip�Q۳Q���}�x�JvTZ�_A�RY��o@REDsUC�S�FIT���PRJвQ�l2LI�NE_XYSKIp.sM���5VIAF7� � @HDt�s �$JO ���$Z_UPLy ��ZT���m�����_M�i�EP��#�) ��m�=�D�YDЦ�(c��� 5*�P�A5 �CACH�S���p8�@�P�CC��MI�SF���d�T��c֤�$H�Oo@�B!�COM	MMc��O���͗I`g�A�{єPVP�r ��Ѡ��S��ZUp�ذ����4AMP�F�AI��Go�2�A9DA�lRMREДa���GP�
p���S�YNBUFvVVR�TD��䠱OL�E_2D_q3��W.63PC_v`Us�yQG���ECCU�x�VEM�p��b�VIRCA�ś�ҟ�_DELA�s�A� �� �dAG��RqXYb��CqW�qs���F��1 �T`rIM�Y��;�@ W�GRA�BB1Y.s3�LE�R<pC���F_D�`��+&50������R ջ��7P��LASs���_GEĥ� �@��A$��TT���Aa,P6" uI{�r?�BG�_LEVEat`PaKtpA��A͗GID NO,Qq�qA O�n�Я�"O�Sc�.�N$�T�LAŤ��R�C�ױ`'#��D�!DE� ��A:�P:�dp�CAT <��@�2�T A �-$5#�iNQ%Dq!Ȥ�o T��ؑnd@� $#AIT�"�<��eSh�SFaPƣ�  � 'k^�fpUR�� SM�%s��"�HADJ��u��ZD�� D���AL��`��л��PERI��$MoSG_Q�$�ю�AC�4B�d@�����!M������W)N�`�D� �ܡ�M�`�q �"`C��`0$�"�0�BJ�4s���Qpb@&6WN��P�XVR�C��,�T_OVR~'�ZABC_E���rg2���
����X!ACTVS�� � � $�5<1q"CTIV屭��IOmb�3���QITlcprDVP
pq��@�`,��A�0P	S���B Z��B�Ѡp�1��LST�R�ѱ�l�1E_S�Q<�X!DCSCH�B� L�SD�5O�P���P����GNp$Ds<��S@_FUN����6�ZI�%��	g�$L����pZMPCFk5�"�@6��A�aLNK�
��Ak�l4� �$��}�4CMCMD���SC_Q.Q�P�1? $JLSFTD��RRcR\W hU `FWπքaR�WUX~�5UXE)q�V~�WU �UmU�Q�Q�Y�Q�WKP�FTF?�RSd��Z�%��"<(�D�%"&aYM�D�� g� 8f�հIU)3�HEIGH\s�?(��&����&`��� � �灅0�$B�t�uq�SH�IF��<(RV��F ���b\0C��GR<Q 0��Gr�aPS���YDx�CE0V���C%aSPHERE�� ,�ahwo�i��$��# 1 �����q���ДA @	� @@3#���s�r�v��w~�v�
]b�so�@��q �q8��� ���q��� 1�}T�uB���0\�t���_��q�N�BANFWD � �s�q��K ^ݰ1 1�u߀��04EOA�T w/o pasrt_���	� �r4��%�j�I�[��� ���֟��ǟ���� �!�3�E�W�i�{���Hү��ɇ2Ԍ�q4��  �<��ݰA3����1�ɇ4N�`�r���ɇ5����ſ׿ɇ6����*�ɇA7G�Y�k�}�ɇ8��0�Ͼ���ɇMA��& ά�  ���OV_LD  ���0��Ʉ�`�! ׋r�`HѼߎ�U@?� M��
���!����UP�D��p�H�<�F�ɂ_�C� �! �p�'q��X���CHKf������rz�c�u�RSS����q������C@���y_GӀ��
 4���A�F�w� j��������������� =0B���"�2�d�M���� ������� #�F�>]b� ��}�������<��V 1�u��>�q�[�l��%0G_IN�0�qd���dO&MASS\/ �Zp'MN[/�#MO�N_QUEUE ��u��@�@*�N]�U��N�&�(��#END�!��)EaX@?�#@BE0��/�#�c�'�� eqR�AM %�*%�� /���"TASKhqN?��O A�/xrߵ?�0DATA�s]�;@�v2�u WOiO{O�O�OJO�O�O �O�O_�O/_A_S_e_^OINFO�s5M��$!_�_�_�_�_o o*o<oNo`oro�o�o �o�o�o�o�o&4�W�T	5L P	�1~~�DIT 
�?����4WERFL�-8B#��RGADJ7 uzA�Π�t�?� �uc!�v�!�0}C��?���9z#&EA<@�R�V�%�T��xP�/A2Y�Ur	H� l#'yA"�>���Хw�t$Ć*Ӏ=/Ղ **:ނ� �я����u����С��qC�R=� �s��-�[�Q�c�ݟ ����ǟ��ϟI��� 3�)�;���_�q����� ��!�˯ݯ����� 7�I�w�m�������� �ٿ�e��!�O�E� W���{ύϻϱ���=� ����'��/ߩ�S�e� �߉ߛ��������� ��+�=�k�a�s��� ���������Y��� C�9�K���o������� ��1����#�@GY�}�:&	O (� O:ŉqǃ�=�9���PR�EF �� �� 
)$RIORI�TY�'�&��qMP�DSPk1�z�R/'U��'���vODUCT��1�zE169511��0���_TG�p�2yzn"HIBIT_DO-?�l$TOENT 1�u{ (!AF_INEY ?7?!tcp??=�!ud.?g>!icmV?]�n"kXY
�u|�Q�)� ��?�?	 ��?O�5�?2OOVO =OOO�OsO�O�O�O�O �O
_�O._@_*m#
����RB��_�_<�>W�����/��@r_�_���Qm�u�A3�?,  � [q@0oBoTofo�u���V�Z�_�o�o�o�o�S�USENHANCE� a]_rAwkdx�_<#u  �j&��|& .v1�qPOR_T_NUMZ#	 ��%�q_CAR�TREP� �<"S�KSTAY'�+SL�GS	0�;���SUnothingD%�7�I�Y���|���������pT?EMP })����m�_a_seiban���,� R�=�v�a��������� �͟ߟ��<�'�`� K���o�������ޯɯ ��&��J�5�G��� k�����ȿ���׿�� "��F�1�j�Uώ�y� �ϝϯ��������0� �T�?�dߊ�u߮ߙ���߽������,�  �$H ���sVE�RSI8 {'}� �disabl�eVp��SAVE �}*	267_0H705/����!,����h?� !	5�c"�g�^��S�e{���������������ro��_�  �1�;�� �}'I�l~�^�URGE�`B� �.�1WF� �!\$}b��&W0�D!�zWR�UP_DELAY� �}@&�_HOT %}%e"+�O�R_NORM�AL.�">�bS�EMIr��L!Q/SKIPJlw[x�/�@/R/d/'- Q�/�/�/�/�/�/? �/?7?I?[?!??m? �?�?�?�?�?�?�?!O 3OEOOiOWOyO�O�O �O�O�O�O__/_�O�?_e_S_�_�_�_]�RACFG ��l;���Q_PA�RAM�3�; Dzh@`�d�2Cp�;�@�}pCv�qBBH>�RBTIF�~�PCVTMOU�w��u��PDCR�J� ��3!?�ͦB?�"Bɳ@�5�?�8�;s彰'-�����Y�?����Sq*/�&.;e�m2r��KZ;�=g;�?4�<<�� 8p�} �� ������%�7��I�[�m��RDIO�_TYPE  �Qaw�EDPRO[T_�Q �B��0[a�EL`Ň�2�!Ջ �^qB� X`�*�^P�t�_� ����+�ɟ��{/� o_!�#�5�k�Y���}� ����ߟ�ie����� 1��U�C�e�g�y��� ѯֿ�������-�� Q�?�u�cϙϻ���߿ ���ύ���;�)�K� q�_ߕ߷ϼ��ϝ�w� ����7�%�[�I�� �ߦ��w���s����� ��!�W�E�{���� ����������� A/Q�����kcŇ?INT 2"1�=��aG;� ���;�[��f�0  4FcfWvx� �����//>/ ,/b/H/Z/�/�/�/�/ �/�/�/??:?(?^? p?V?�?�?�?�?�?�? �?O O6O$OFOlORO�O~O�O�^EFPO�S1 1#�� @ x�Y�c	 +__O_[X�O_A_�_ �_�_a_�_�_o�_o Do�_hoo�o'o�o�o ]ooo�o
�o.�oR �ovs�G�k ���*����r� ]���1���U�ޏy�ۏ ���8�ӏ\������� -�?�y�ڟş����"� ��F��C�|����;� į_���������B� -�f����%���I��� ��ϣ�,�ǿP�b� ���IϪϕ���i��� ��߱��L���p�� ��/߸���e�w߱�� ��6���Z���~��{� ��O���s���� �2� �����z�e���9��� ]���������@�� d����5G�� ��*�N�K ��C�g�/ ���J/5/n/	/�/ -/�/Q/�/�/�/?�/ 4?�/X?j???Q?�? �?�?q?�?�?O�?O TO�?xOO�O7O�O�O mOO�O__>_�Ob_ �O�_!_�_�_W_�_{_ o�_(o:o�_�_!o�o mo�oAo�oeo�o�o�o $�oH�ol�� =O�����2� �V��S���'���K� ԏo���
������R� =�v����5���Y��� �������<�ן`�r� ��Y�����ޯy�� ��&���#�\������ ��?�ȿڿu�����"� �F��j�ώ�)ϋ� ��_��σ�ߧ�0�B� ����)ߊ�u߮�I��� m��ߑ���,���P��� t����E�W���� �����:���^���[� ��/���S���w�  ������ZE~� =�a��� � D�hz'a� ���
/�./�+/ d/��/#/�/G/�/�/��$REFPOS�2 1$����1 @ x}/�/�/G?2?k? q/�?*?�?N?�?�?�? O�?1O�?UOgOOO NO�O�O�OnO�O�O_ �O_Q_�Ou__�_4_ �_�_j_|_�_oo;o �__o�_�oo�o�oTo �oxo�o%7�o�o j�>�b� ��!��E��i�� ����:�L����ҏ� ��/�ʏS��P���$� ��H�џl�������� �O�:�s����2��� V���񯌯���9�ԯ ]�o�
��V�����ۿ v�����#Ͼ� �Y��� }�ϡ�<�����rτ� ���
�C���g�ߋ� &߈���\��߀�	�� -�?�����&��r�� F���j������)��� M���q������B�T� ��������7��[ ��X�,�P�t ����WB{ �:�^��� /�A/�e/w//$/ ^/�/�/�/~/?�/+? �/(?a?�/�? ?�?D? �?�?z?�?�?'OOKO �?oO
O�O.O�O�OdO �O�O_�O5_G_�O�O ._�_z_�_N_�_r_�_ �_�_1o�_Uo�_yoo �o�oJo\o�o�o�o �o?�oc�o`�4 �X�|���� �_�J������B�ˏ f�ȏ���%���I�� m���,�f�ǟ��� �����3�Ο0�i�� ��(���L�կ篂��� ί/��S��w���� 6���ѿl�����ϴ� =�O����6ϗςϻ� V���z�ߞ� �9��� ]��ρ�ߥ߷�R�d� ������#��G���k� �h��<���`���� �������g�R��� &���J���n���	�� -��Q��u�"4�n��� �$R�EFPOS3 1�%��� @ x� ��dO���G �k�/�*/�N/ �r/�//1/k/�/�/ �/�/?�/8?�/5?n? 	?�?-?�?Q?�?�?�? �?�?4OOXO�?|OO �O;O�O�OqO�O�O_ �OB_T_�O_;_�_�_ �_[_�__o�_o>o �_bo�_�o!o�o�oWo io�o�o(�oL�o pm�A�e� ��$����l�W� ��+���O�؏s�Տ� ��2�͏V��z���'� 9�s�ԟ��������� @�۟=�v����5��� Y��������ۯ<�'� `��������C���޿ y�ϝ�&���J�\��� 	�CϤϏ���c��χ� ߫��F���j�ߎ� )߲���_�q߫���� 0���T���x��u�� I���m�����,��� ���t�_���3���W� ��{�����:��^ ����/A{��  �$�H�E~ �=�a��� ��D///h//�/'/ �/K/�/�/�/
?�/.? �/R?d?�/?K?�?�? �?k?�?�?O�?ONO �?rOO�O1O�O�OgO yO�O_�O8_�O\_�O �__}_�_Q_�_u_�_ �_"o4o�_�_o|ogo �o;o�o_o�o�o�o �oB�of��7 I�����,�� P��M���!���E�Ώ i��������L�7� p����/���S���� �����6�џZ�l�� �S�����دs�����  ����V��z���� 9�¿Կo������� @�ۿd�����#υϾ� Y���}�ߡ�*�<��� ��#߄�oߨ�C���g� �ߋ���&���J���n� 	���?�Q����������$REFP�OS4 1&����;� @ x������� l�������d������� #��G��k�� <N����1 �U�R�&�J �n�	/���Q/ </u//�/4/�/X/�/ �/�/?�/;?�/_?q? ??X?�?�?�?x?O �?%O�?"O[O�?OO �O>O�O�OtO�O�O!_ _E_�Oi__�_(_�_ �_^_�_�_o�_/oAo �_�_(o�oto�oHo�o lo�o�o�o+�oO�o s��DV�� ���9��]��Z� ��.���R�ۏv���� ������Y�D�}���� <�ş`�������� C�ޟg�y��&�`��� ��寀�	���-�ȯ*� c�����"���F�Ͽ� |���ȿ)��M��q� ϕ�0ϒ���f��ϊ� ߮�7�I�����0ߑ� |ߵ�P���t��ߘ��� 3���W���{���� L�^���������A� ��e� �b���6���Z� ��~����� a L� �D�h� �'�K�o� .h����/ �5/�2/k//�/*/ �/N/�/�/�/�/�/1? ?U?�/y??�?8?�? �?n?�?�?O�??OQO �?�?8O�O�O�OXO�O |O_�O_;_�O__�O �__�_�_T_f_�_o �_%o�_Io�_moojo �o>o�obo�o�o! �o�oiT�(� L�p���/�� S��w���$�6�p�я ���������=�؏:� s����2���V�ߟ� ����؟9�$�]����� ���@���ۯv����� #���G�Y����@��� ��ſ`�鿄�Ϩ�
� C�޿g�ϋ�&ϯ��π\�nϨ�	���-�:���$REFPOS5 1'���X�� @ x���� ߞ߉����� �߁�
���@���d� �߈�#���Y�k�� ���*���N���r�� o���C���g����� &����nY�- �Q�u��4 �X�|�);u ����/�B/� ?/x//�/7/�/[/�/ �/�/�/�/>?)?b?�/ �?!?�?E?�?�?{?O �?(O�?LO^O�?OEO �O�O�OeO�O�O_�O _H_�Ol__�_+_�_ �_a_s_�_o�_2o�_ Vo�_zoowo�oKo�o oo�o�o.�o�o va�5�Y�} ���<��`���� ��1�C�}�ޏɏ��� &���J��G������ ?�ȟc��������� F�1�j����)���M� ��诃����0�˯T� f���M�����ҿm� ����ϵ��P��t� Ϙ�3ϼ���i�{ϵ� ��:���^��ς�� ߸�S���w� ��$� 6������~�i��=� ��a������ ���D� ��h������9�K��� ����
��.��R�� O�#�G�k� ���N9r �1�U���/ �8/�\/n/	//U/ �/�/�/u/�/�/"?�/ ?X?�/|??�?;?�? �?q?�?�?O	OBO�? fOO�O%O�O�O[O�O O_�O,_>_�O�O%_ �_q_�_E_�_i_�_�_ �_(o�_Lo�_poo�o �oAoSo�o�o�o�o 6�oZ�oW�+� O�s����� V�A�z����9�]� ���������@�ۏd� v��#�]������}� ���*�ş'�`����� ���C�̯ޯy���ů�&��J�W��$RE�FPOS6 1(����u�? @ x�� =�����߿�Ϟ�'� ¿$�]�����ϥ�@� ����vψ���#��G� ��k�ߏ�*ߌ���`� �߄���1�C����� *��v��J���n��� ����-���Q���u�� ����F�X������� ��;��_��\�0 �T�x�� �[F�>� b���!/�E/� i/{//(/b/�/�/�/ �/?�//?�/,?e? ? �?$?�?H?�?�?~?�? �?+OOOO�?sOO�O 2O�O�OhO�O�O_�O 9_K_�O�O2_�_~_�_ R_�_v_�_�_�_5o�_ Yo�_}oo�o�oNo`o �o�o�o�oC�og d�8�\�� 	�����c�N��� "���F�Ϗj�̏��� )�ďM��q����0� j�˟������7� ҟ4�m����,���P� ٯ믆���ү3��W� �{����:���տp� ����ϸ�A�S�� � :ϛφϿ�Z���~�� ���=���a��υ� � �߻�V�hߢ����'� ��K���o�
�l��@� ��d�����#����� 
�k�V���*���N��� r�����1��U�� y�&8r��� ��?�<u �4�X���� �;/&/_/��//�/ B/�/�/x/?�/%?�/ I?[?�/?B?�?�?�? b?�?�?O�?OEO�? iOO�O(O�O�O^OpO �O_�O/_�OS_�Ow_ _t_�_H_�_l_�_�_ o+o�_�_oso^o�o 2o�oVo�ozo�o�o 9�o]�o��.@ z����#��G� �D�}����<�ŏ`� ��������C�.�g��t��$REFPO�S7 1)������ @ x� �Z�؟ß ��� ���D�ߟA�z� ���9�¯]������ ��߯@�+�d�����#� ��G����}�ϡ�*� ſN�`����GϨϓ� ��g��ϋ�߯��J� ��n�	ߒ�-߶���c� u߯����4���X��� |��y��M���q��� ���0������x�c� ��7���[������ ��>��b����3 E���(� L�I��A� e� /���H/3/ l//�/+/�/O/�/�/ �/?�/2?�/V?h?? ?O?�?�?�?o?�?�? O�?ORO�?vOO�O 5O�O�OkO}O�O__ <_�O`_�O�__�_�_ U_�_y_o�_&o8o�_ �_o�oko�o?o�oco �o�o�o"�oF�oj ��;M��� ��0��T��Q��� %���I�ҏm������ ���P�;�t����3� ��W���򟍟���:� ՟^�p���W����� ܯw� ���$���!�Z� ��~����=�ƿؿs� ���� ��D�߿h�� ��'ω���]��ρ�
� ��.�@�����'߈�s� ��G���k��ߏ���*� ��N���r����C� U���������8��� \���Y���-���Q��� u���������XC |�;�_�� ��B�fx %_���/� ,/�)/b/��/!/�/ E/�/�/{/�/�/(?? L?�/p??�?/?�?�? e?�?�?O�?6OHO�? �?/O�O{O�OOO�OsO �O�O�O2_�OV_�Oz_ _�_�_K_]_�_�_�_ o�_@o�_do�_ao�o 5o�oYo�o}o�o��o�o`K��y�$�REFPOS8 �1*����q� @ x +=w���=� �a��^���2���V� ߏz�������]� H������@�ɟd�Ɵ ����#���G��k�}� �*�d�ů��鯄�� ��1�̯.�g����&� ��J�ӿ忀���̿-� �Q��u�ϙ�4ϖ� ��j��ώ�߲�;�M� ����4ߕ߀߹�T��� x�����7���[��� ����P�b���� ��!���E���i��f� ��:���^����� ����eP�$� H�l��+� O�s� 2l� ���/�9/�6/ o/
/�/./�/R/�/�/ �/�/�/5? ?Y?�/}? ?�?<?�?�?r?�?�? O�?COUO�?O<O�O �O�O\O�O�O	_�O_ ?_�Oc_�O�_"_�_�_ X_j_�_o�_)o�_Mo �_qoono�oBo�ofo �o�o%�o�om X�,�P�t� ��3��W��{��� (�:�t�Տ������� ��A�܏>�w����6� ��Z��������ܟ=� (�a����� ���D��� ߯z����'�¯K�]� ��
�D�����ɿd�� ��Ϭ��G��k�� ��*ϳ���`�rϬ�� ��1���U���y��v� ��J���n��ߒ��-� �����u�`��4�� X���|������;��� _������0�B�|��� ����%��I��F �>�b�� ���E0i� (�L���/� //�S/e/ //L/�/ �/�/l/�/�/?�/? O?�/s??�?2?�?�? h?z?�?O O9O�?]O �?�OO~O�ORO�OvO �O�O#_5_�O�O_}_�h_�_�Y�$REF�POSMASK �1+����Q� �R@��_�W�WXNO  ��_�_�^MOTE�  l�TEa_CFOG ,LmgQ>T��b�QPL_RAN�GHaBQe��fOW_ER -e�`��fSM_DRYP�RG %i�%�I_�o�eTART �.�nzUME_�PRO�o�oc�T_�EXEC_ENB�  �e�iGSP�D<p~p�x�xT3DB��zRM��x�INGVERSI_ON jR��YI_AIRPUR�` DzdY��[�MIeb/LnBR� ��` ;)y�MOVH`������P<Ō�mz�~q �2m  >T\fT!� >W��@�R�d�v�|� X�b4��PC3ґ�����@��H�A�;f�`˷�@��[�]�������@�ᾲ�}g���@���!� d�_��_/��$� e� ���D��������s�T_�PT�`Jk�e�OBOT_ISOLCl�Ԡա�e�U^�NAME
���~A�_CATEGh��cc`������O�RD_NUM ?��hR�H?705  >T������PPC_TI�MEOUT�o x��PS232eb13�e�s LT�EACH PEN�DAN/�aW����؍H_FPMai�ntenance Cons��|�>U�"��BTNo Use؏�Ϗ������8#�5�D�NPOp1®�a�cD�C7H_L?p4	�С�	�с�!UD�1:�߃�R�PVA�IḺ1×��e�D�PACE1 2=5k�߀jW܏��d�b��ի���< �U�?� ����������,� M�\�T�f�x��<��� ��������1F gb�t�������\�� ���@�Q8f �����j� /��>/_/6/t/�/ ������/�/ (?I?�/�/?f?�?�? �/�/�/�/�?
??6O @?OlO�OdOvO�O�? �?�?�?O�O*OLOV_ w_6_�O�_�_�_�_�O �O__&_8_J_l_vo Do�o�o�o�o�o�_ o"o4o�oXozo�� d����� 0BT�x���� ȏ�����.�,�>� P�b��������ӟ�� �	���?�:�L�^� p���4���ȟү��� �)��>�_�Z�l�~� ��B�����a���� 7��L�m�h�z����� ��b�Կ�� �!���j� W�>�lߍ߈ϚϬϾ� p���������D�e� <�N�w�ߨߺ����� ���$�.�O����� l��������������� �"�D�Nr�� |��������� 0R\}<��� ����,� Pr|/��/�/�/�/ �////(/:/�/^/ �/�?�?j?�?�?�?�? O?$?6?H?Z?O~? �?�O�?zO�O_�O_ 7_2ODOVOhO_�O�O �_9_�_�_o�_$oEo @_R_d_v_�_:o�_�_ �o�o�oBo/De `oro�o�oH�o�o� �o��=��&�O�n ����h���� '��p�]�D�r����� ����ď֏����&� ��J�k�}�T�f����� ��ҟ䟖��*�4�U� �j���r�������ί �����(�J�TϚ� xϙϫϒϔ�޿ܿ�  ����6�X�b߃�B� �߹ߠ����������  �2���V�x߂���R���������� ��$RSPACE2 25���0�� ��0�B���f�� ����������<�3-�?�Q�c�u�' �����F�98NoMCE4bt ���\� /{��M/n/E/�/�/�CE5������/ /5/L?�/,?�?�?z?8�?�?�/CE6�/�/ �/??�?8?j?�O�?�aO�O�O�O�O_�?CE7OO%O7OIO�O mO�O�__�_�_o�_8"oCo!_CE86_H_ Z_l_~_0o�_�_�oOo��o!BWxVoC�EG 9nk� �jt
�p �  ne���"� 4�F�X�pc�hw��op��t֏��d��� �#�5�G�Y�k�}�s� ������şכ����� �9�K�]�o������� ����������� ��Y�k�}���������໯ͯ߯�� `S @LŴ�Z�6�>���µ#ϩϻ� ���ʜ����"�@��� (�j�|�F�P�bߔ��� �ߪ߼���0�B�`�� H���f�p�����Ƽ
z�K�s�Y_MODE  nk�a�S :ni� :����ovϟ����
	:b�TMgP mf�`�o o�o���o�o����0Ef�|CWORK_ADq����*��!R  ��{`�?�_INTVALq������OPTI�ON� ��!V�_DATA_GR�P 2≮��D2�P'G/#k/V) $��/�/�/�/�/�/? �/??(?^?L?�?p? �?�?�?�?�? O�?$O OHO6OlOZO|O~O�O �O�O�O�O_�O2_ _ B_h_V_�_z_�_�_�_ �_�_�_�_.ooRo@o vodo�o�o�o�o�o�o �o<*LN` ����������8�&�\�t��$S�AF_DO_PULSq�u�l��v�CAN_TIMp��B����R =�#h�#�{~�]%]
��a!]�~ց3� `/� �2� D�V�h���������Xԟ�t#l��2�ց�d�*�\"ԃ�O��st�І�Z>���P���B�_ @T�  T���������T D��B�T�f�x� ��������ҿ���� �,�>�P�b�_��P�r�r��υ��  �;��oV��~p��
�u��Di|�S  � �� ~ޅ΁��^�p߂� �ߦ߸������� �� $�6�H�Z�l�~��� ����������� �2� D�V�h�z���������@������
V�m� J\n����� �)��*<N `r������0k�4�+�ۈ����� ////A/S/e/w/�/ �/�/�/�/�/�/?? +?=?O?a?s?�?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O 4�O�O_#_5_G_Y_ k_}_�_��_�_�_�_��_oo1oCo�4�M�DЀo`jao`o`�����o�o�o�o �o�g�o�o"4F Xj|����� ����0�B�T�f� x���������ҏ���@��,�>�P�%��y� )�[�������Ο��� ��(�:�L�^�p���������ƪ��ϯ��.����������	123456�78K�h!BQ!��'Z�����l�~����� ��ƿؿ������%� 7�I�[�m�ϑϣϵ� ���������!�3�E� V��yߋߝ߯����� ����	��-�?�Q�c� u���X�j������� ��)�;�M�_�q��� �������������� %7I[m�� �����!3 Ei{���� ���////A/S/ e/w/�/�/Z�/�/�/ �/??+?=?O?a?s? �?�?�?�?�?�?�?�/ O'O9OKO]OoO�O�O �O�O�O�O�O�O_#_ 5_G_Ok_}_�_�_�_ �_�_�_�_oo1oCo@Uogoyo�o�o<�i� �o�o�eb_�o	o�Cz  A�a�_   �s�2��}Q�jׇ <�
sw�/  	�<�2�o������|psa��l� �*�<�N�`�r����� ����̏ޏ����&�@8�J�\�n����(up��(������ϟ�� ��)�;�M�_�q��� ������˯ݯ����<��a�qYr<7�� -��q  �G�a�Ksy�D��q>�qt  Np��0��tp���� `3rD��п�A}y��6�3r��$SCR_GRP� 1?#�`�#��� 	$ ��`r Tu	 �D�� L�]�V��o͑�iǗ�8�Ͼ�*}�cp��?D1� D�~c��׻��
CRX�-10iA/L �23456789�0�p2� @уp�2�L O�3q
V?14.00 lЌȴR�z�s{ ��@L���;���;��)�bq[ɏ���	�������� �2�B����H�L���P���G�5_�B�m�D�%�C6&�C�3���5��B��sh�C3ґ�����@��^�A�;}�`˿�@��NB�  =�8B�ovD%�C6 �L��3q�����#�0w��i/xh7p,��B�  B�n�l��rh�ANp��  @6p̬�h�@���� ?	���h�Hr�����h�F@ F�` �;&_Jo� ����`�����0�)B�7� }h������ �/
/C/./g/y/� �çϙ'�/q�
�/�/��@-;��6p0?r��F71=�V7Uv�b��?51��&�5 ���3��0��23q �2�3�1�?OM�1(H4OFOO��|O�O@�?�/�O�O�O��0߀f4�3!W�O>_���ECLVL  3qg���ҷ0j7\Q�L_DEFAUL�TdTW����6pxSHOTS�TR�]�1�RMIP_OWERFcP2ux�U[R�PWFDO�V� �ZRVENT� 1@kQkQ�S �L!DUM_E�IPJ_���j!?AF_INE�PIo���!FToxnD?o�o!;´o�L��o��o!RPC_MAI���I��o4�c'VIS�I�#�?!OPCU41�摗o�!TMP�pPU�2id���!
PMON_�PROXY�5fe �d��r2�.mfS����!RDM_SR�V��2ig����!�Rh4�3hh�H�!%
�`M{�/li7����!RLSYNC̕���8����!gROSo��4ϟ�,�!
CE�pMT'COM-�5fk�x�{!	A�CONSy��4glg�į!A�WOASRCˏ5fm��v�!A�USB��3hn��\�!STM�Pv�1joK����o�̿����L_�QICE�_KL ?%k� (%SVCPGRG1��=�'�2=�DB�,�3e�j�,�4��D��,�5�Ϻ�,�6����,�7�
�,�]�M�H�9U�Z�)���� ,�/Ϫ�,�W���,�� ��,���"�,���J�,� ��r�,�ߚ�,�G��� ,�o���T����T��� :�T���b�T���T� 8��T�`���T��� T���*T���RT� � z|�(����,��%� �
��2VA ze������ �//@/+/d/O/v/ �/�/�/�/�/�/?�/ *?<?'?`?K?�?o?�? �?�?�?�?O�?&OO JO5OnOYO�O�O�O�O �O�O�O_�O4__F_�j_U_�_ �_DEV� i�U�T1:���4~�TGRP 2De��P!�bx 	_� 
 ,�P�Q �_o�T.o@o'odoKo �o�o�o�o�o�o�o�o �o<#`rY� }{�U���yo�� $��H�/�l�~�e��� ��Ə؏����� �2� �V��z���C���� C�ܟß ����6�� Z�A�S���w�����د �ѯ�e���D���h� O�������¿����� ߿��@�R�9�v�]� �ρϓ���'���߽� *��N�5�G߄�kߨ� �����������&�8� �\�C����϶�m� ���������4�F�-� j�Q���u��������� ��B��7x /������� ,P7t�m �����/[(/ :/!/^/E/�/i/{/�/ �/�/�/ ??�/6?? Z?l?S?�?w?�?�?/ �?�?O OODO+OhO zOaO�O�O�O�O�O�O �O__@_R_9_v_�Y�d �Xzh96�T 	 A���:�A�36|=>���h�@�- �Z��P�G�A=���?�&%�H��@�������]B���A|������?����§=������]@��}����AÖ@���h����A�Z��Y%PR�OVA�_Xo���la�Qle|o�gto��o�o�o�o�o y%�Yo'  �o�oJ �n���
�. �"��2�4�F�|�j� ���Ǐ������� �.�0�B�x�����ޏ h�ҟ�������*� ����w���P�����ί �����X�=�|�� p��������ʿ��� 0��T�޿H�6�l�Z� |Ϣϐ������,϶�  ��D�2�h�V�xߞ� ����ߎ������
� @�.�d�ߋ��T�v� P��������<�~� c���,����������� ����V�;z�n \������. R�F4jX� |���*�/ /B/0/f/T/�/��/ �z/�/v/�/??>? ,?b?�/�?�/R?�?�? �?�?�?OO:O|?aO �?*O�O�O�O�O�O�O �O_TO9_xO_l_Z_ �_~_�_�_�__�_o �_�_�_2ohoVo�ozo �o�_�oo�o
�o .dR��o��o x������*� `�����P�����ޏ ̏����h���_��� 8���������ڟȟ�� @�%�d��X��h��� |�����֯���<�Ư 0��T�B�d���x��� �տ������,�� P�>�`φ�ȿ���v� �������(��Lߎ� s߅�<�^�8ߦ�����  ���$�f�K���~� l����������>� #�b���V�D�z�h��� ���������:���. R@vd��� ���*N <r���b�^ �/�&//J/�q/ �:/�/�/�/�/�/�/ �/"?d/I?�/?|?j? �?�?�?�?�?�?<?!O `?�?TOBOxOfO�O�O �OO�O�O�O�O�O_ P_>_t_b_�_�O�_�O �_�_�_oooLo:o po�_�o�_`o�o�o�o �o�o H�oo�o 8������� PvG�� �z�h��� �����(��L�֏ @�ҏP�v�d�������  ��$�����<�*� L�r�`���؟������ �ޯ��8�&�H�n� ����ԯ^�ȿ���ڿ ���4�v�[�m�$�F�  ώ��ϲ������N� 3�r���f�T�v�xߊ� �߮���&��J���>� ,�b�P�r�t����� ��"����:�(�^� L�n����������� �� 6$Z��� ��J�F��� �2tY�"�z �����
/L1/ p�d/R/�/v/�/�/ �/�/$/	?H/�/<?*? `?N?�?r?�?�/�?�? �?�?�?O8O&O\OJO �O�?�O�?pO�O�O�O �O�O4_"_X_�O_�O H_�_�_�_�_�_�_�_ 0or_Wo�_ o�oxo�o �o�o�o�o8o^o/no bP�t��� �4�(��8�^� L���p����͏���  ��$��4�Z�H�~� �����n�؟Ɵ���  ��0�V���}���F� ����ԯ¯����^� C�U��.��v����� п����6��Z��N� <�^�`�rϨϖ���� ��2ϼ�&��J�8�Z� \�nߤ�����
ߔ��� ��"��F�4�V���� ����|���������� �B���i���2���.� ����������\�A ��
tb���� ��4X�L: p^����� 0�$//H/6/l/Z/ �/��/�/�/�/|/�/  ??D?2?h?�/�?�/ X?�?�?�?�?�?O
O @O�?gO�?0O�O�O�O �O�O�O�O_ZO?_~O _r_`_�_�_�_�_�_  _F_oV_�_Jo8ono \o�o�o�o�_�oo�o �o F4jX� �o��o~���� �B�0�f�����V� �����ҏ����>� ��e���.��������� ��Ο�F�+�=���� �^���������ܯ� �B�̯6�$�F�H�Z� ��~�����ۿ���� ��2� �B�D�Vό�ο ���|�����
���.� �>ߔϺϋ���d߾� ���������*�l�Q� ���������� ���D�)�h���\�J� ��n���������� @���4"XF|j ������� 0TBx��� h�d�/�,// P/�w/�@/�/�/�/ �/�/?�/(?j/O?�/ ?�?p?�?�?�?�?�?  OB?'Of?�?ZOHO~O lO�O�O�OO.O�O>O �O2_ _V_D_z_h_�_ �O�__�_�_�_o.o oRo@ovo�_�o�_fo �o�o�o�o*N �ou�o>���� �� �&�hM��u�p��$SERV_MAIL  �u�����ql�OUT�PUTw���p@l�RV 2�E�i��  (��R�ޏl�SAVE�����TOP10 �2F�� d 76�� (�F� X�j�|�������ğ֟ �����0�B�T�f� x���������ү��� ��,�>�P�b�t��� ������ο���Ϙ(�:��YP����F�ZN_CFG G����t����r�GRP 2H�|�	� ,B  � A���qD;� �B���  B4~�sRB21�oHELLu�I���ˀ̏��%�4�%RSR4�5�G߀� kߤߏ��߳������� "��F�1�j�U���~���  �h��%����������	�b�p����ބw
��2�pd�	������HK 1J�� "������������� ��61CU~y���������OMM K��5���FTOV_ENB�w�h��HOW_R�EG_UIU��IMIOFWDL �L$�ŊWAIT�R��²��vܿ��TIMv����VAv���_�UNITQ &�L]CoTRYv��l�MB_HDD�N 2M��  ����u� ��/��/ �/�/�/�/"??+?X?^2r!Eu�N�ɧ�Y�tp3��O|; �����<�u>(z5���X�p��<,��?�  �?�;�Ʉ� _�" k 9�pG�y:`4@nv�=�=@�v���JE�tG@��`G�MON_AL�IAS ?e$ǀhe=��O�O�O�O �J�O__/_A_�Oe_ w_�_�_�_X_�_�_�_ oo�_=oOoaoso�o 0o�o�o�o�o�o�o '9K�oo��� �b����#�� G�Y�k�}���:���ŏ ׏鏔���1�C�U�  �y���������l�� ��	��-�؟Q�c�u� ��2�����ϯ�󯞯 �)�;�M�_�
����� ����˿v����%� 7��[�m�ϑ�<ϵ� �������Ϩ�!�3�E� W�i�ߍߟ߱����� ������/���@�e� w���F�������� ���+�=�O�a�s�� ������������ '9��]o��� P�����5 GYk}(��� ���//1/C/� g/y/�/�/�/Z/�/�/ �/	??�/??Q?c?u? �?2?�?�?�?�?�?O O)O;OMO�?qO�O�O��O�ObC�$SMO�N_DEFPRO�G &�����A &�*SYSTEM*��O�O�BRECAL�L ?}�I ( �}kOO_a_s_�_�_�_ =_�_�_�_o o(o�_Lo^opo�o�o �o9o�o�o�o $ �oHZl~��5 ����� ��D� V�h�z�����1�ԏ ���
����@�R�d� v�����-���П��� ��*���N�`�r��� ����;�̯ޯ��� &���J�\�n������� 7�ȿڿ����"ϵ� F�X�j�|ώϠ�3��� �������߱�B�T� f�xߊߜ�/������� �����+�P�b�t� ����=�������� �(���L�^�p����� ��9������� $ ��HZl~��5 ���� �D Vhz��1�� ��
//�@/R/d/ v/�/�/-/�/�/�/�/ ??*?�/N?`?r?�? �?�?;?�?�?�?OO &O�?JO\OnO�O�O�O 7O�O�O�O�O_"_�O F_X_j_|_�_�_3_�_ �_�_�_oo�_BoTo foxo�o�o/o�o�o�o �o�o+Pbt ���=���� �(��L�^�p����� ��9�ʏ܏� ��$�����$SNPX_�ASG 2P����J��� P 0 '�%R[1]@1�.1+���?���% u���M���ȟ{����� �"����X�;�M���⸀u�����abX ��诛�ݯ�q�B��� 7�x�+�m�����ҿ� ǿ����>���b�E�@WϘ�[����ϸ�&� �Ϫ���-߀�Q��F� ��:�|߽ߠ������� ����M���q�T�f���jߜ��︁�4 �������>���b�� W���K��������� ��(^���e w�{����� H�=~1�U ����/A2/D/ '/h/�]/�/�/�/� �/�/�/�/.??R?5? G?�?k?}?�?�/�?�?�?O��OGOJ/<O }O�?�O�?�O�O�O�O _�O1__&_g_J_\_��_�_�_�_�_�_�X% �_'oZOo]o@o�o�_ o�o�O�o�o�o�oGʨn�7x+ m����~����ko�>�!�=�PAR�AM QJ�^T� �	��P�e글����� ���=�OFT_K�B_CFG  ��tQ�:�OPIN_�SIM  J���������[�RV�NORDY_DO�  ��ǅ/�QSTP_DSBێ���s�Wx[�SR �Rމ � &���OS2  OR�T�Wy�u��TM_CTL 3Sޅ���  p% |�	��-���B�Q�[t ��|���1�C�^sށ_� �������˯�^� p��%�7�I�ʿܿ� ������6�H�Z�������GRPۈ�p����OP_ON_E�RR<���PTN ��D��RING_PRM���N�VCNT_GP� 2Tޅ����x 	��`�_pN߇�r�̫ߊ�VD5Т�1Uj����і������� 
��.�U�R�d�v�� ������������ *�<�N�`�r������� ��������&8 J\n����� ���"4Fm j|������ �/3/0/B/T/f/x/ �/�/�/�/�/�/�/? ?,?>?P?b?t?�?�? �?�?�?�?�?OO(O :OLO^O�O�O�O�O�O �O�O�O __$_K_H_ Z_l_~_�_�_�_�_�_ �_oo o2oDoVoho zo�o�o�o�o�o�o�o 
.@Rdv� �������� *�<�c�`�r������������PRG_CO+UN��͔����'ENB��M����_UPD 1V>��T  
Ϗ&� b�t���������Ο�� ���?�:�L�^��� ������ϯʯܯ�� �$�6�_�Z�l�~��� ����ƿ�����7� 2�D�V��zόϞ��� �������
��.�W� R�d�vߟߚ߬߾��� �����/�*�<�N�w� r���������� ��&�O�J�\�n��� ��������������' "4Foj|��������،_INFO 1WP��6�X	 �<3��?��?��>^.�D=P`;������/�^v?���?�Z�>�\�F=#�;�czC3ґ���Փ@��A���5�`�?@��&z�=�@ �>/ȝ ����CD2MD�4��Ca����'��N&/�8'�YSDEBU)G��Q��%d�a SP_PASS���B?s+LOG �XMZ�  z%�!?���%�,  �5�%UD1:\�$3�"o_MPC�/ �$(�",?�,�(2�/2?SAV Y�)��؉�!(:�(SV�`;TEM_TIM�E 1Z�'[�� 0  Q��-�2?�3�3MEM�BK  P�5��� �/5OGOWLX�|6�� @WO$��yO�O�LrO�O,�Jn! �@�1_ (_:_L_�3d_v_�_�_�_�_�_ ��_�_o o,o>oPoboto�o��e�o�o�o�o�o &8J\n�����������5S!K@H�� K �_��q�eGM�`T�L�  D�O�� ��5�A�O���O�H	A�_��E�W�%`Q_��  ���H�M�lȟڟ ߏ ����B��7�I�[�m��%U�����o˯!{ӯ��	��-�?� Q�c�u���������Ͽ�����)�9T1SVGUNSP����# 's%�D�2�MODE_LIMG [�9w"@�2M��m�\�-?�ABU�I_DCS _3�s!#@�������C 2������C *���=� 
C�,=�@��W�(�7X��,��EDIT `����&9�  E�;���CZ  C�$H��SCRN �a�-���0��-,)� �cD��	0OG b���؅6����SK_OPTI�ONh Iw!��_D�I� ENB  ��s%��BC2_G_RP 2d���� X�ϺD�PC8����a?%�����CFI��f��&=��(?C� o�������������� �� 9$IoZ �~������ �5 YD}h� �������/+/ =/�a/L/q/�/�/�/ ��3��/@� �/?�/ (??L?:?p?^?�?�? �?�?�?�?�?O O6O $OFOlOZO�O~O�O�O �O�O�O�O�O2_X�� F_X_v_�_�__�_�_ �_�_�_o*o<o
o`o No�oro�o�o�o�o�o �o&J8n\ ~������� � �"�4�j�X���D_ ����֏���x��� .�T�B�x�����j��� ���ҟ�����,� b�P���t�����ί�� ޯ��(��L�:�p� ^�������ʿ��� ��6�H�Z�ؿ~�l� �ϴϢ��������� � �D�2�h�V�x�zߌ� �߰�����
���.�� >�d�R��v����� ��������*��N�� f�x�������8����� ��8J\*� n������� "F4jX�| �����/�0/ /@/B/T/�/x/�/d� �/�/�/??�/>?,? N?t?b?�?�?�?�?�? �?O�?(OO8O:OLO �OpO�O�O�O�O�O�O �O$__H_6_l_Z_�_ ~_�_�_�_�_�_o�/ &o8oVohozo�_�o�o �o�o�o�o
�o@ .dR�v��� ����*��N�<� ^���r�����̏���� ޏ ���J�8�n�$o ������ȟڟX������4�"�X�B�v��$�TBCSG_GR�P 2gB���  �v� 
 ?�  �� ����ׯ�������1���U�g�z���i��_d�H��?v�	 HA���e��>���>f���\e�AT��A ���пܸ�����G��?L��Ʋpܿ޾�;ff�������v�򾺠$�l�@��R����ff>�33��e�~�B˿m��J�����Ɍ�϶�҃�H��B����B��϶�K�E�K�j�}� H�Zߨ��ߐߢ�������ؐ6�	V3�.00��	cr;xl�	*X�P�u���[���H���� q��p��  O��Cp�����z�J2ʁ�k�����#�	 @����8�J�\�n��������������CFoG mB���Y ��#����9#�/�/U (���s���� ��*N9r ]������� /�8/#/\/G/�/�/ }/�/�/�/�/�/?3 ��?.?@?�/s?^?�? �?�?�?�?�?�?O'O 9OKOOoOZO�O~O�O �Ov�b��O>��O __ H_6_l_Z_�_~_�_�_ �_�_�_o�_2o oVo Dofohozo�o�o�o�o �o�o
,R@v d�������� ��<�*�`�N���r� ����̏ޏ������ 8�&�\�n�����L��� ��ڟȟ����4�"� X�F�|�j�������֯ į�����B�0�R� T�f����������ҿ ����>��V�h�z� $ϪϘϺϼ������ (��L�^�p߂�@ߦ� ���߸��� ��$��� 4�Z�H�~�l����� �������� ��D�2� h�V���z��������� ��
��.>@R �v������� ��N<r`� �����//� $/J/8/n/\/�/�/�/ �/�/�/�/?�/ ?F? 4?j?X?�?|?�?�?�? �?�?O�?0OOTOBO xOfO�O�O�O�O�O�O �O__*_,_>_t_� �_�_�_Z_�_�_�_o o:o(o^oLo�o�o�o �ovo�o�o �o6 HZ&�~�� �����2� �V� D�z�h��������� ����
�@�.�d�R� t����������П� ��_0�B��_����r� ����̯��ܯ��&� 8�J�����n����� ȿڿ�����"��2� 4�F�|�jϠώ��ϲ� ��������B�0�f� Tߊ�xߚߜ߮����� ���,��P�>�`�� t��$�V������� ��L�:�p�^����� ���������� " $6l~��\� ���� 2 hV�z���� �
/�.//R/@/v/ d/�/�/�/�/�/�/�/ ??<?N?��f?x?�? 4?�?�?�?�?�?�?O 8O&O\OnO�O�OPO�O�O�O�O�O�N  $P(S (V<_(R��$TBJOP_�GRP 2n�E��  �?���C(R	�TR[Spb\��@��X  �(U�P �, � ��P^(S @$P?�Q	 �A����U?C�  DBW�Q��Q>tP>\?�`�UaG�:��o�];ߴAgT���U�QA�:c��UKoVg�_�_>�Q��\)?���f8�Q��Q�RL��>y�.`$P;iG,b��gAp:`�`Do�oA�ff�eto�T�`xr'~:VM�,b���`Qt<om(U@�;�R�uCр�Q��Q�u�t�b�e�ff��u:�6/�q?�{33�uB   �q �����r�a�d�}^<�:�S��~��px}�����@��H���$��x-q�p�u=�`<�#�
(v�QtP;/��ڨ�?��P�B�
��%�0i�U0�fw X�B�P�~�����D�Ο �ҟ���?��ԟ^��x�b�p���ϯ(SC��(V���U	V3�.00yScrxl�T*��T#Q��at3� F�� H�H F6�� F^ F��� F�f F�� G� G5� G<
 G^]� G� G����G�*�G�S� G�; G���C�Dup��E[�� E� F(� F-� FU`� F}  F�N� F� F��� Fͺ F�� F�V G�� Gz Ga� 9ѷ챸�HD �d�2_�*�(V�.� ��U��F^ED_TCH qb[�)�0�
(  ��u$Pd$%�����(TB�����C��U���STPARS  �X��TPHR �A�BLE 1rbYC L����C� �0#�������'W/Q*��	��
����Zժ(Q������N7�RDIB�lQY�@k�}ߏߡ߳��O#�5�?�Q�c�u��;�S!�jS ��H�Z�l�~� ��������������  2DVhz�� G] �$�kRX��	���� ����߼���������;��NUM  V�ElQ�P0P� W��;�_CFGG s�[�Q@TP�IMEBF_TT�&�V����VER��Q&�R 1=tJ� 8��(R�#Pc! �@�   K/]/o/�/�/�/�/�/ �/�/�/?#?5?G?Y? k?}?�?�?�?�?O�?��?OO1OCN� WOiOCN!S�O�O�O�O �O�O�O_"_4_F_X_ j_|_�_�_�_�_�_�_ �_oo0oBoTofj0$�_�&@'%��L�IF u���"!��d"!�d(�D�
����@pd� d	}��`SC�RN v� �IOx_CUR ew����	)D��O{PREV �xc}�VtS��2y�c{ xDO��) ��}g1���m�b�l�d��qMI_CH�AN� '% e�D_BGLVL����e�ETHERADW ?*����.��0Ā:eǀ4:�7d:bc:db� ďc׏dd�d�e��ROUT !��!�8�w�h�?SNMASK��'#~��255.v���t��������OOLOFS_DI&��՚�ORQCTRL zJۓ�/��T�:�L�^�p��� ������ʯܯ� �� $�6�H�Z�j����|����}�PE_DET�AI��ۚPGL_�CONFIG ������/c�ell/$CID?$/grp1��+� =�O�a�sώ���� ���������χ��.� @�R�d�v�ߚ߬߾� �����߃ߕ�*�<�N� `�r��������� �����&�8�J�\�n� ���!������������}��FXj|@��s������� �!3EW��{ �����d�/ ///A/S/e/��/�/ �/�/�/�/r/??+? =?O?a?�/�?�?�?�? �?�?�?�?O'O9OKO ]OoO�?�O�O�O�O�O �O|O_#_5_G_Y_k_ }__�_�_�_�_�_�_ �_o1oCoUogoyoo �o�o�o�o�o�o	���User �View �}}�1234567890:L^p����t ��� y2 -y�o��"�4�F�X���'r3�����ʏ@܏� �_�!��~4�� Z�l�~��������՟�~5I�� �2�D�V�h�ǟ���~6��¯ԯ����
��{�=��~7 ��v���������п/���~8e�*�<�N�`��rτ�㿥ϫ� �lCamera+z!������ �2�D�"E��n߀ߒ�8��߾����������  ���y��V�h�z�� ���W�������C��@.�@�R�d�v������ �����������
 ��@Rd����� �������H�y. @Rdv�/�� ��//*/</N/ ���"���/�/�/�/ �/�/�?,?>?�/b? t?�?�?�?�?c/�Ű� Q?OO*O<ONO`O? �O�O�O�?�O�O�O_ _&_�?��d��Or_�_ �_�_�_�_sO�_oo __8oJo\ono�o�o9_ ���)o�o�o& 8�_\n��o��@�����o�g9� ?�Q�c�u�����@�� ϏᏈ��)�;�M�(_�q� �	��0���� ��П������*�<� N���r���������̯ s�������p�%�7�I� [�m��&�����ǿ� ����!�3�E���� 9�ܿ�ϣϵ������� ���!�3�~�W�i�{� �ߟ߱�Xϒ���H��� �!�3�E�W���{�� �������������� ������i�{����� ����j�����V�/ ASew�0���}+  ���/�� Sew����� ������;�A/S/ e/w/�/�/B�/�/�/ ./??+?=?O?a?-  )�?�?�? �?�?�?�?O O2ODOVK   f?}Oh? VOx:�O�O�O�O__ )_;_M___q_�_�_�_ �_�_�_�_oo%o7o Io[omoo�o�o�o�o �o�o�o!3EW i{������A}
 (  �0( 	 ��� 2� �V�D�z�h��������ԏ�����J�J ̰/a�s��� �/����͟ߟ��
# P�-�?�Q���u����� ����ϯ����^� ;�M�_�q�����ܯ�� ˿ݿ$���%�7�I� [Ϣ����ϣϵ����� �����!�3�z�W�i� {��ϟ߱��������� @��/�A��e�w�� ���������� `�=�O�a�s������� ������&�'9 K]�������� ���#j|Y k}������ �B/1/C/�g/y/ �/�/�/�//�/�/	? P/-???Q?c?u?�?�/ �/�?�?�?(?OO)O ;OMO_O�?�O�O�O�? �O�O�O__%_lOI_ [_m_�O�_�_�_�_�_8�_2_�@ bo�,o>ocg�p���"frh:\tp�gl\robot�s\crxxa10�ia_l.xml �_�o�o�o�o�o�o0+=O��Pu �������� �)�;�RL�q����� ����ˏݏ���%� 7�N�H�m�������� ǟٟ����!�3�J� D�i�{�������ïկ �����/�F�@�e� w���������ѿ��� ��+�B�<�a�sυ� �ϩϻ��������� '�>�8�]�o߁ߓߥ� �����������#�5�:Wh�Q ob`�<< `` ?�5�x�5�p����� �������,��$�F� t�Z�|����������������(6V<P(��$TPGL_OUTPUT �@Q�@QS   h}������ �1CUgy �������	/�/hX��- cel�l/floor/�wall 8901234567P/ b/t/�/�/�%6R- �/ �/�/�/??�/�/J?@\?n?�?�?�?<7}�? �?�?�?	OO�?�?QO cOuO�O�O�OCO�O�O �O__)_�O7___q_ �_�_�_?_Q_�_�_o o%o7o�_Eomoo�o �o�oMo�o�o�o! 3�o�oi{��� �[����/�A� �O�w���������W� i�����+�=�O�� ]���������͟e�۟���'�9�K��2 $$%/�� ������ׯɯ���� �C�5�g�Y���}��� ��ӿſ�����?�@1�c�Uχ�yϫ�}S�����������0�@�Z�T�f�`� ( 	 �ϛ߉߿߭� ���������+�a� O��s�������� ���'��K�9�o�]�������������3&�  <<�� "4m [mG� �-*���� �Rd�h�4 ����//v / N/�:/�/�/p/�/�/ */�/??�/8?J?$? V?�?�/�/�?�?b?�? �?�?�?4OFO�?jO|O OhO�O�O�O�O�OXO _0_�O_f_x_R_�_ �__�_�_�_�_o,o o4obo�_Jo�o�oDo �o�o�o�oto�oL ^�oj�n��� :����H�Z�4� ~����x�Ə`����� ��2�D���,�z��� &�����Ο��V�h� .�@�ڟH�v�P�b��� ���������*����`�r�)WG?L1.XML0ߧ���$TPOFF_�LIM 	 =�����N_S]V��  7�Ϻ�P_MON ��Ѵ=�=�2���STRTCHK' �϶�ϸ��VTCOMPAT��n�ӶVWVAR� ����� KE� ��=�����_DEFPR�OG %3�%�ROS�߱�_DISPLAYİ�3���INST_M�SK  +� ~�INUSERd���LCKm�4�QU?ICKMEN���oSCRE��~o�tpscԠm�����ϲ��_��S�Tb�ϹRACE_�CFG ������	��
?�~,�HNL 2�����P�� ������������.�I�TEM 2�p�� �%$1234?567890W�i�  =<a�������  !������ k�����U�y�9K ��a�����	�- ���u���� 7����)�M _q��A/g/y/� �///%/�/�/[/? -?�/9?�/�/�?�/�? ?�?�?E?�?i?�?DO �?_O�?oO�O�OO�O /OAOSO�OwO#_I_[_ �O_�O�O_�_�_=_ �_os_o�_�_ro�_ �o�_�o�o'o�oKo]o &�oA�oQw�o�o �o+5�Y�+� =��a����c�� ��ߏ�U���y����� !�o�ӏ����	���-� ?��c�#���G�Y��� o��3����ׯ;�� ����+�����˯E� ﯛ���ӿ7���[�m� ��ϵ�uχ�뿓� �!���E��i�)�;�@��Q����Ϟ�*�S6���<���  ��� H�����
� �-��Q����UD1:\^������R_GRP 1��D�� 	 @@������������#���3�J�X���^��m�����?�  ���������� ;)KM_�� �����7�	q�K]��SC�B 2���  �������//�'/9/��UTORIAL ���E�/���V_CONFIG ���C���A���/�-OUTPUT� ���� ���/3?E?W?i?{?�? �?�?�?�?�?�?O�!  ?3OEOWOiO{O�O�O �O�O�O�O�O_O/_ A_S_e_w_�_�_�_�_ �_�_�_o_+o=oOo aoso�o�o�o�o�o�o �o&o9K]o �������� �"5�G�Y�k�}��� ����ŏ׏����� 1�C�U�g�y������� ��ӟ���	��,�?� Q�c�u���������ϯ ����(�;�M�_� q���������˿ݿ� ��$�7�I�[�m�� �ϣϵ���������� !߽/�%?_�q߃ߕ� �߹���������%� 7�*�[�m����� ���������!�3�D� W�i�{����������� ����/AR�e w������� +=Nas� ������// '/9/J]/o/�/�/�/ �/�/�/�/�/?#?5? G?X/k?}?�?�?�?�? �?�?�?OO1OCOT? gOyO�O�O�O�O�O�O �O	__-_?_POc_u_ �_�_�_�_�_�_�_o o)o;oMo^_qo�o�o �o�o�o�o�o%�7I,���� hzdqS�H��� ���#�5�G�Y�k� }�����Toŏ׏��� ��1�C�U�g�y��� ������ӟ���	�� -�?�Q�c�u������� ��ϯ����)�;� M�_�q���������˿ ݿ���%�7�I�[� m�ϑϣϵ�ƿ���� ���!�3�E�W�i�{� �ߟ߱���������� �/�A�S�e�w��� �����������+� =�O�a�s��������� ������'9K ]o������� ��#5GYk�}�����$T�X_SCREEN� 1�|u�dp�}ipn�l/�gen.htm�/'/9/K/]/�� Panel� setupa,}�/pip/rm�i_log.txta/�/�/�/�/�/q �RMI_LOG�/ }�?>?P?b?t?�?�?,?"?�?�? �?OO)O�?MO�?qO �O�O�O�O�OBOTO_ _%_7_I_[_�O _�O �_�_�_�_�_�_t_!o �_EoWoio{o�o�oo (o�o�o�o/�o �o�ow������H��UALRM_MSG ?��� ��
*�<� m�`�����������؏�ޏ��3�&�W��S�EV  ����	�ECFG ���  ��@�  A�� �  B��
  X�������"�4� F�X�j�|����������GRP 2���� 0�	 ?��1�>��q�(�P���i��?� ��^�I_BB�L_NOTE ����T��#l�������DEFPR0?%� (%K�r�� �`�����ROS2 ��x�ƿ�ֿ���3���W�B�{ύ��FK�EYDATA 1y���p ��� ������6�0�� �2��,(��c���Qߎ�u�ANCE�L����}�REV �STEP����EX�T���{�INIS�H�F�}�ORE INFOG�J��� �������������;�M�4�q�X������ ��/frh�/gui/whi�tehome.png������
.�/Sew����<FRH/FCG�TP/wzcancel����!<3�prev�m����Dwznext\�//'/�9/�wzfinish�w/�/�/�/�/N-infof/�/	? ?-???:c?u?�?�? �?�?L?�?�?OO)O ;OMO�?qO�O�O�O�O �OZO�O__%_7_I_ �Om__�_�_�_�_�_ h_�_o!o3oEoWo�_ {o�o�o�o�o�o���o /ASelo� �����r�� +�=�O�a��s����� ��͏ߏ񏀏�'�9� K�]�o���������ɟ ۟�|���#�5�G�Y� k�}������ůׯ� �����1�C�U�g�y� �������ӿ���	� ��-�?�Q�c�uχ�� �Ͻ�������ߔ�� ;�M�_�q߃ߕ�$߹�@��������� ���������I�[�m�E���{�, ����������,�� P�7�t���m������� ������(:!^ E�i�����  �o6HZl~ ��ߴ����/  /�D/V/h/z/�/�/ -/�/�/�/�/
??�/ @?R?d?v?�?�?�?;? �?�?�?OO*O�?NO `OrO�O�O�O7O�O�O �O__&_8_�O\_n_ �_�_�_�_E_�_�_�_ o"o4o�_Xojo|o�o �o�o�oSo�o�o 0B�ofx��� �O����,�>� P�'t���������Ώ ����(�:�L�^� 폂�������ʟܟk�  ��$�6�H�Z��~� ������Ưد�y��  �2�D�V�h������� ��¿Կ�u�
��.� @�R�d�v�ϚϬϾ� �����σ��*�<�N� `�r�ߖߨߺ����� ����&�8�J�\�n� ������������� ��"�4�F�X�j�|����e����e����������������,�B�fM �������� >P7t[� ������/(/ /L/3/p/�/a��/�/ �/�/�/ ?�$?6?H? Z?l?~?�??�?�?�? �?�?O�?2ODOVOhO zO�OO�O�O�O�O�O 
__�O@_R_d_v_�_ �_)_�_�_�_�_oo �_<oNo`oro�o�o�o 7o�o�o�o&�o J\n���3� ����"�4��X� j�|�������A�֏� ����0���T�f�x� ���������/���� �,�>�E�b�t����� ����ί]����(� :�L�ۯp��������� ʿY�� ��$�6�H� Z��~ϐϢϴ����� g���� �2�D�V��� zߌߞ߰�������u� 
��.�@�R�d��߈� ��������q��� *�<�N�`�r������ ���������&8 J\n����������Ր �>Ր���); M%o�[,m/� e/���/�0// T/f/M/�/q/�/�/�/ �/�/???>?%?b? I?�?�??�?�?�?�? џO(O:OLO^OpO �O�O�O�O�O�O _�O $_6_H_Z_l_~__�_ �_�_�_�_�_�_ o2o DoVohozo�oo�o�o �o�o�o
�o.@R dv����� ����<�N�`�r� ����%���̏ޏ��� ���8�J�\�n����� ��3�ȟڟ����"� ��F�X�j�|�����/� į֯�����0�O T�f�x���������ҿ �����,�>�Ϳb� tφϘϪϼ�K����� ��(�:���^�p߂� �ߦ߸���Y��� �� $�6�H���l�~��� ����U������ �2� D�V���z��������� ��c���
.@R ��v������ q*<N`� ������m/�/&/8/J/\/n/E��p+�E�����/�/�-�/�/�/�&,�?"?�?F?-?j?|? c?�?�?�?�?�?�?�? O0OOTO;OxO�OqO �O�O�O�O�O_�O,_ _P_b_A��_�_�_�_ �_�_�oo(o:oLo ^opo�_�o�o�o�o�o �o}o$6HZl �o������� � �2�D�V�h�z�	� ����ԏ������ .�@�R�d�v������ ��П������*�<� N�`�r��������̯ ޯ�����8�J�\� n�����!���ȿڿ� ��ϟ�4�F�X�j�|� �Ϡ�w_��������� �%�B�T�f�xߊߜ� ��=���������,� ��P�b�t����9� ��������(�:��� ^�p���������G��� �� $6��Zl ~����U��  2D�hz� ���Q��
// ./@/R/�v/�/�/�/ �/�/_/�/??*?<? N?�/r?�?�?�?�?�?��?���;������	OO-MOOOaO;F,M_�OE_�O �O�O�O�O_�O4_F_ -_j_Q_�_�_�_�_�_ �_�_�_ooBo)ofo xo_o�o�o�o�o���o ,>P_?t� �����o�� (�:�L�^�������� ��ʏ܏k� ��$�6� H�Z�l���������Ɵ ؟�y�� �2�D�V� h���������¯ԯ� �����.�@�R�d�v� �������п����� �*�<�N�`�rτ�� �Ϻ�������ߑ�&� 8�J�\�n߀�ߤ߶� ����������o4�F� X�j�|��߲����� ��������B�T�f� x�����+��������� ��>Pbt� ��9��� (�L^p��� 5��� //$/6/ �Z/l/~/�/�/�/C/ �/�/�/? ?2?�/V? h?z?�?�?�?�?Q?�? �?
OO.O@O�?dOvO �O�O�O�OMO�O�O_�_*_<_N_%�P[}�%����y_@�_�]u_�_�_�V,�o o�o&ooJo\oCo�o go�o�o�o�o�o�o �o4XjQ�u �������0� B�!�f�x��������� �O�����,�>�P� ߏt���������Ο]� ���(�:�L�۟p� ��������ʯܯk� � �$�6�H�Z��~��� ����ƿؿg���� � 2�D�V�h����Ϟϰ� ������u�
��.�@� R�d��ψߚ߬߾��� ���߃��*�<�N�`� r����������� ��&�8�J�\�n��� W�������������� "4FXj|� ������0 BTfx��� ���//�>/P/ b/t/�/�/'/�/�/�/ �/??�/:?L?^?p? �?�?�?5?�?�?�? O O$O�?HOZOlO~O�O �O1O�O�O�O�O_ _ 2_�OV_h_z_�_�_�_ ?_�_�_�_
oo.o�_ Rodovo�o�o�o�o����k�������o�o}�o/Av,-�r%��}� �����&��J� 1�n���g�����ȏڏ �����"�	�F�X�?� |�c�������֟��� ��0�?oT�f�x��� ������O������ ,�>�ͯb�t������� ��K�����(�:� L�ۿpςϔϦϸ��� Y��� ��$�6�H��� l�~ߐߢߴ�����g� ��� �2�D�V���z� ��������c���
� �.�@�R�d������ ��������q�* <N`������ ���ǟ&8J \nu����� ���"/4/F/X/j/ |//�/�/�/�/�/�/ �/?0?B?T?f?x?�? ?�?�?�?�?�?O�? ,O>OPObOtO�OO�O �O�O�O�O__�O:_ L_^_p_�_�_#_�_�_ �_�_ oo�_6oHoZo lo~o�o�o1o�o�o�o �o �oDVhz ��-����
�h�.�0�����Y�k�}�U�������,��⏕� ��*�<�#�`�G��� ��}�����ޟ�ן� ��8�J�1�n�U���y� ��ȯ���ӯ�"� F�X�j�|������Ŀ ֿ�����0Ͽ�T� f�xϊϜϮ�=����� ����,߻�P�b�t� �ߘߪ߼�K������ �(�:���^�p��� ���G����� ��$� 6�H���l�~������� ��U����� 2D ��hz����� c�
.@R� v�����_� //*/</N/`/7��/ �/�/�/�/�/�?? &?8?J?\?n?�/�?�? �?�?�?�?{?O"O4O FOXOjO�?�O�O�O�O �O�O�O�O_0_B_T_ f_x__�_�_�_�_�_ �_�_o,o>oPoboto �oo�o�o�o�o�o �o(:L^p� ����� ��� 6�H�Z�l�~������ Ə؏������2�D��V�h�z������$U�I_INUSER  �������  �����_MENH�IST 1����  (� ̐��'/S�OFTPART/�GENLINK?�current=�menupage�,71,1 15 ޟS�e�w��)�*�1��=�ůׯ�������37=��Z�l��~��* �2�8<�16��߿�ϒ�����ȱ30�c�uχ��(�:�3ï�������Ϲ�7�4��f�xߊ�0��#�=�ö22������$���*��7�B�T�f�x����  >�������	��-��� Q�c�u�������:��� ����);��_ q����H�� %7�[m ����V��/ !/3/E/0�i/{/�/�/ �/�/�/��/??/? A?S?�/w?�?�?�?�? �?`?�?OO+O=OOO aO�?�O�O�O�O�O�O nO__'_9_K_]_�O �_�_�_�_�_�_�_|_ o#o5oGoYokoV/to �o�o�o�o�o�o�_ 1CUgy�� ������-�?� Q�c�u��������Ϗ �����)�;�M�_� q��������˟ݟ� ����7�I�[�m�� ��|o*�ǯٯ���� !�$�E�W�i�{����� .�ÿտ�����/� ��S�e�wωϛϭ�<� ��������+ߺ�O� a�s߅ߗߩ߻�J��� ����'�9���]�o�������$U�I_PANEDA�TA 1�������  �	�}3htt�p://1.1.�0.10:308�0/frh/jc�gtp/flex�dev.stm?�_width=0�  _dummy.htm��K�]���)pri9�����}������������ )7[B �x�������3E,i�����  � r������ �� /S$/��H/Z/ l/~/�/�/	/�/�/�/ �/�/ ?2??V?=?z? �?s?�?�?�?�?�?
O} ��)E��E/JO\O nO�O�O�O�?�O;/�O �O_"_4_F_�Oj_|_ c_�_�_�_�_�_�_�_ ooBoTo;oxo_o�o �o!O3O�o�o, >�ob�O���� ���Y��:�!� ^�p�W���{���ʏ�� �Տ�$��H��o�o ~�������Ɵ؟+��� ��2�D�V�h�z��� 󟰯��ԯ�ͯ
�� .�@�'�d�K������� �����U�g�%�*�<� N�`�rτ�׿����� ������&ߍ�J�\� C߀�gߤ߶ߝ����� ����"�4��X�?�|� ������������� �q�B���f�x����� ������9����� >P7t[��� ����(��� ^p����� �a�/$/6/H/Z/l/ ��/w/�/�/�/�/�/ ? ??D?+?h?z?a?`�?�?�?5G}��?@OO0OBOTOfO)�? �O�zO�O�O�O�O�O _xO5__Y_@_R_�_ v_�_�_�_�_�_o�_�1oCo*ogo�QK��$UI_POST�YPE  Q�� 	 �so�o�bQUICK�MEN  �k��o�o�`RESTO�RE 1�Q�  ��*defaul�t�SING�LE}PRI�Mmmenu�page,74,1t����u� ��,�>�P��t��� ������OuZoя�U� �0�B�T�f�x���� ����ҟ䟇���,� >�P���]�o���󟼯 ί�����(�:�L� ^�p���%�����ʿܿ ����ϑ�Z�l� ~ϐϢ�E��������� ߱�2�D�V�h�z�%� /ߙ߫������
�� .�@���d�v����O����������mS�CRE�`?�m�u1sc9p�u2Y�3Y�4Y�5*Y�6Y�7Y�8Y�6�wTAT�m� �c<Q�jUSER;�@��R�ks[���3��4���5��6��7��8���`NDO_CFG ��k�0�1�`�OP_CRM5 c �5=�`PD������No�ne�b��_INF�O 2�Q� �`0%$����� �BT7x [������/��l�OFFSET' ��i�/�� 2p��Y/k/}/�/�/�/ �/�/�/�/E/�/L?C? U?�?y?�?�?�?�?�? ;�oMOBO
2OgO���I�WORK �� OVO�O�O|/��UFRAM]p�V�RTOL_A�BRT_�REN�B'_XGRP 1��-y�aCz  A�}S{Q��{_�_�_�_�_�V�_�_Z�`�UGX[6[MSK � JU�6[NQ�%�	�%�?�o8U_'EVN&PJd<�fv.3�7+
 h[�UEV&P!�td:\event_user\�oF�`C7�oDO[ FtM��`SP�a�gsp�otweld}!C6W%7[�zd!zo�o���w2a� ��$�Y�����:� ��^�p��������ʏ ܏�g�V���6�H�~� ӟ������-�؟Q� c�� ���D���h�z���fW�@3���SA8��!�3� �X�j� E�����{�Ŀֿ���� ��0�B��f�x�S� �Ϯω����Ͽ�����,��$VARS__CONFI1 �7+� FP���3�C�MRcR2�7+�+i[ 	\ �B%�1: SC130EF2 *�߼п䥙�8�{�2`�S  �[?��P@�Pp:�P�-� �O���;�M�z��uﴢ���UA�������� B����������f� C��g�R���v����� ����<���Q��u�;�GRID6�b�O� �?���}p�>L���@��?� ?,g?��33��  @��@��>��.P������?�IA�D��M~�,		��eWeG�P ��xyH>�ISIO�NTMOU�o �����b8�c�rQ �FR:\�\DA�TA�   �wUD1�LOG�7  �EX����' B@ ��@"��^/�v/��/�� � n?6  �����=!�,g�'5�  =�����!��� -TR�AIN'/�!�"�rd3p�%�(7#KT�t�{ҭ�k (> (9x=6	x?�?�?�?�? �?�?O OO$O6OHO�ZOlO9�IS_GE����k�`.P��
wP.P�B�G$ RE� �jY��;�LEX��D�� 1-e��VMPHASE'  �e���>��RTD_FILT�ER 2��k �����_�_�_�_ �_�_�_o#o5o��~_ couo�o�o�o�o�o�o��o�	SHIFTMENU 1�[;/
 <M,%M/c���Ag�w� �������T��+�=���a�s������	LIVE/SN�A_�%vsflsiv&^ҏ��� SETU_���menu����o����R!u��[9�wM�O��^�z=�Z%D����O��<0�@��$WAITDINEND�D1��	�OK  ��$��r?�SS�&�TIM���~�G���2��ëR���q�����$�RELE=Qӧ��	��<��_ACT�Ҩt:$�_� �2��%��ӿ8և�RD�IS_�T�	�NSP��왴��{��3��r�<#��1:�XVRQ��^�$ZABCvz�1�� ,0
AD02ۿ�⑌�VSPT ��\��$
n�n����N� �߽�DCSCH��2E0�
�A y�I����@�����߹�MPC�F_G 1�<�0@��$�6���ÿ��ZE1p���>�D018
����Q`� �G����<?����=�?�\��?�ʿ��|>��I��.J����CD2LD4��D0�0�A@H����V=��O>��ă�{q=�y�0���G�٣���?�O��x����s����}+��l�.L���}���zD4�������T�=�����}��=�Q��� |�g���>�������Ca���?�+��N��*��������P��q���� )7 a����1�57�I��u��P����_C_YLINDcQ��� �& ,(  *&7##`G�k ���� � /p%///[/ �/�/�/��/b/H/ �/�/!??v/W?i?���2���� � �?4ݗ��?��ONh�?AOז[AA���SPHERE 2�̻/�O?�O�O �O�O9?LO'_9_�/]_ �O�O�_z_�_�__�_ �_F_X_5o�_Yo@oRo��o�_�o�o�oy�ZZq� ǰ�