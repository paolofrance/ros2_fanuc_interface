��  ��A��*SYST�EM*��V9.4�0341 1/�17/2024 A�  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  ��4�ADV_I�N� 0  0KO�PEN� CRO �%$CLOS\� %EDI�BA �"IO_CNV�� l� RAC��LO�MOD_wTYP@FIR��HAL�#IN_;OU�FAC� g�INTERCEP:fB: SIZ@!�LRM_RECO�N"  � ALM��"=!  �&ON\�!� MDG/ �$DEBUG1PA2d43AO� �o"��!_IF�� � $ENA�BL@�#� P dj�#UU5K51MA�h� 2�
� OG�|f Z0CURR_�1:P $�3LIN@�1:�4$�$AUSO[4�� OD/2$SEV�_AND_NOA��2TP8"�6�4�5��APPINFOE=Q/  �L ��0�1EA H �GD9EQUI�P 38@NA�M/0�\B_OV�R�$VERS�I� �!PCOU�PLEm  	 �$�!PP�1CESI0�2�G101"P�0�B
 � $�SOFT�T_I�D�3OTAL_E%Q00�1�@N" �@U SPI
 �0^�E�X�3CRE ]Dn�BSIGz@�O|�K�@PK_FII0�	$THKY�RWPANE�D ~� DUMMY1d�yT!1�U4�Q���AR�1R� � $TITI1� ��0�Td�T!0��T�P�T5�V6�V7
�V8�V9�W �U�W@Q�U�W�Q�U�W1�WU1�W1g1g2b~�SBN_CF�![6@$L!J� �; K2A_CMNT��$FLAGS�]�CHE["$�b_OPTzB � �ELLSETUP�  `8@HO,h@I PR�1%�c#�	qREPRx�0D�+�@�+r{3uHM�I MN<% UTO�BZ U�0� D9DEVIC&�STI_@�� �@�r3�dpB�d�"VA�L3ISP_UN9I��p_DO�v7�yFR_FP�%�1�3��A`s�C_W�A�t\q�OFF_��@N�DEL1�L��0�q�1<��r?�q=�SS?��`2QRU1��#Z�;QTB1��b�MO� 1�E "REM1�����wREV�BILǇ��!XI� ��R 7 � OD�`끿$NO�`M@�������/�"���� �/��PD��d p E R�D_E〘�$F�SSB+6�`KBD�_SE�uAG� G
#Ba"_��2��� �VQ�{5�`X��C  %�`q_8"�@2�rD�$!S�]D6 P�A�Q#�B;���_�OKa��0m P_C�� ��`t�U pLACI�!q>���� ��qCOMM� # $D:�P�P=�ٙz_��R'@BIGALL;OW� (K�2:]BPVAR���!�	Q�#BL�@� �C ,K�qΤ�`S���@M_O]�����CCFS_UTӀ@�"�AS�'-��[pXw��b@ 4�0IMCM0�3S@�p�i�ʀi H�_D��<$ G��MA� hT�IMPEE_F�������� ���ǳD_�ӵ÷�DθF��4�_8H��@ T8@|��|�DI��@w�H�� =�PA�C$I?�W�M��F�d7 X8@GR�@�z�M��NFLI�<�ü@UIRE�y4<$2� SWIT~$p0k_N�`S02CF�0�M�,C@S��D��!�Ħ`-�<�J�`J�tV%�k E���.�p p(ڗELBOF� �IշI�p@p0���3�0��� F�2����BA��r�1J1,��z _T!��3p���g3p��rxPVCz� D��CLLB�`P=$�����F��G�� ��0WARNM�p��HK�`���`\ � COR-�r�FLTR��TRA�TI T? � $A�CC�qm�0r�r�$ORI�o&��ReT��Sl���HG�0I��T���A�I��T�t��� � &3�aa�N�HDR�2�2�2!J; HS'�!�3"� �$�5"�6"�7"�8"�9��
��
 /B� @0TRQB7�$�f���A����c_Ul���PCO�c  <0�ϒϤ�xE3nB��LLECΒ}!"MULTI�4��"��2QK2M�CHI�LD^�@!��O�@T�M� "W�STY I29r��=��)2������_�c# |@�0E6$�0�¦�`��!�6uTO �E�	EXT����2B2"��_��$�@�	N�p&��ak� %2k�p% q�r���s��^oA&W���A���M���I )% ]TR>� ' L8@{�e#I r<�A��$J�OBç���IGi ( d��// )'r��#�a�Ǧ�_MOR��) �tT�FL1�:RNGUQ��TBA��P��& ���*p1�(D�#@0��!��0;P�p 5�"�*$������q`1w���rJw�_Rh���C�z<Jz�8�<J��D 1�º9)���"'P��Ɓ�P_?pLҴ+ \8@RORpHF@��sIT
�@NOM��@��,D3s:B!ڲUlPMP�� �0�,�P���0��PI��RA��ќѳC[����
$T���MD3$@T��pUpL���e+�AH�r��T1�JE5A����ÀQ�ƌQ8�ƘQ�CYNT�����PDBGD���-^"ޠPU�$j���������AX)��4�T;AI�sBUF\�[YQ�. ���jV�`[PI��-�@P�WEM�XM�Y\P�VF�WSIMQSTO
��$KEE8cPA��є �BRR�C+R��P���/�`��MARqGA��2{�FAC����LEW�1G!�0���(�:����C�$0W���@pJB���?qDEC�jL��e�"����%1 �֐CH�N��MP��$G��@7wt�_PCCU�1g_FPCEPTCbv�v�S��tw�C�П�V0{���q2��JR��/��SEGFR�`IO��!:@ST��LINn��sPV����P]T2 ��rb���r��Ԡ�1�3` +�?��_��2p� ��`��)�j�y��a�SIZ##��t�T`��@�����RS�� .#�s�Ӧypp��pL��
PAp$�CRC��)�CC��&��p�N�bq��br|�MIN@z�bqz1`��4�D�iC��C��	ҕuא�P���� ޘEVޖ:�F*��_�uF��N �<�P�a�ֱh�K�L�A�S2
QVSCA�uPA��ebP��42C{ �SFp4e����r �4P!Ҵ5��	��O�o�g�Ӏ��m��0�VP�b�����Rs�6� @�������e��R@�HANC$LG�O�=��Q$�ND,=���AR�N8�q0ہ����̳ME�ҎИͲ�PǸRA��̳A�Z���
��EO��F�CT�q�`pBB�!S\�`|0ADIm�Om� ��"��!��_�O�O ��#s�G3�!9�BM�P�t��Y&COq�AcES����n�W_���BAS##XYZW�PR ����!�	�gAR_L~ ��7( V�C������KLBB'$g���bшcv�pCEEVр�FORCERQ��+Q'���_AVG�ӱ֫ӇMOMo0���ի�S��TP�����О�i��=���F�d�AYLwOAD�$ER/��t�35B_X�pc1"���QR_FD� 8 Tw`IQ �3e �Ed6:�C�:�MS+`U{
$��p��&)7d���9eRH7EVI��
f�,1o_IDXp$�倀��@�1���&At��@�`R_H�P��: ��3�����W!�� R_��;C �]0��qpM�q��@$PL�A��M��z�!���qF�������_CU�C�20��:��!PL߰���0� ��U5`M
�Um�<nCTITA{
�%_1�qTR �� ={ PAEGED��p�PDT[RE�Md2`AUTH_KEY  ) �A1Dp@J NO�rSZ_��mC>v�
��C߱FNO_HEADE�a�<�E� d�Pph�'��Ut��M�V��md?p�"P��uCIRTR4p4�N��L���C�@��RJ�%�
��Q:�1�@�
B��:�OR!�9�O���M��qUN_O|ðF�$SYS1�P5d�:�X���V�C��pe�DBPXWO�͐ Ap$SK��A�R*�DBT��TkRLBv�AC�p0�D�u���DJ�4� �_���Qm$��y'P5L!��bWA"�� "�cD+Q�'8Q���2>{ UMMY9��"310��PDB��C+"�QPR6�
 ��DKо�D lm��1$;q$��o7�L8E?��ci�@F7?�2�P�CAGV?$��PWENE�@TڢHu?|h3� RECORP2�IH �@L�wD$LK�E$3��R��;�p1��q�_�D���PROS��T�~�W���P0��TR�IG )FPAUS|'C�tETURN'BV�MRX�U��9���0EW��>pSIG�NAL���R$LAxW��E��F$PE�OG$P8��AH�@ƫ�PC�DSi�DO�Iи��2�1c��6GO�_AWAYBMO��q�����!CS��CwSCBۡJ �/q��G��`I�@� �7p��'��6SR@\``ARGAGE��+`��5TlR~�gQKS~�OF�p�KV�0�V_S]�MP�MA2@X_S�$F?RCINI_!U��<�P�$NE�P�V�TLV�ܠK� �z�%RZ�`b��O�2�P�0OVR10��!����$ES�C_p�uDSBI�O�8�`d�©�VIB� �s���e���f��*�SSW.È��VL_���eARM�-��Ra���eSC`�`�T��Q�MP�Ѡrcp�!r4u5O�ESU����sGw�cGw/sGt�s�GtC �Dwɀ'�} O��IqF��qאSB�F�t�G�cgR���7R�v�$VOLT�wN�S�� ��7Q?T������PX�ORQ�F�;���F�DH_THE@�bW��a�^�ALPH^�+������@ F����ɁR M��ӳ��E�p�3a%(2e�1cF�1M�3a!V���Y��Lr˄�INF� �`2bT#HR^ <�h�T԰J�
� V=�!t{!o0��1��2��{��� {�����!�џ��Ӊd d@��ږ��앞��"�� 1П���"�N��؃xCBv�W�INHBM�ILT7@=��d���C �g�T�����aaha�dha`���@Y�AF��O�઩�����ʧ�� a`Nô�稧�R`̩����PL����#���TMOU����C�������c��CA(���?�A�̩��I��B�3DI8����_�STI�ų�۸OX���@����AN���aW$�c������$��	��g�_�����`RA�`�`pfS� ��MCNUa�������VERSP=��_`Ig�F@г�������G�DN"4�G.��ǧ�F�B�Ťק�M�'�F�_�M>ي ���Ýt ��k֝q�dO2 C�`�e������DI� ����#��շ�1҄��g�Fh ���#�O�N�%�a��VAL� �CR��_SIZp��R�+a^�REQ_�R�|�MBR�|�CH a����ʓ��|�����*�^�S_E�vh��gg�FLG���ge$CV�yM7`�a��FLX@�)B#bֵe���5AL�`�C_H��T��W���0�b�s � ��NDMS�'�� ��K.c�`_M@X�STWf� ����AL�`���a����E���E��IAG@�_�to�E�T2	Ap���Q��  �	8p�	Ap�	6�@�_D��!��
�`���6�BpT�� ?�'!Q.�����!L��?`O-Y0P.LD��pS�w!�@�FRI�@ �`����Am��IV!��NA�U�P�`��a��S�L!W����`L-c's'&s�C)g��0 <���1~���d�a�!��w(�����p�"��`�ERSM� P���F@X$ �b�l�tNBAW�q_TB��m�(PNS_PE�A��s�,0���SAV7�(�&WM5��'�CAR��`�1t4��}2CRQ�� 0�d�3qE�P��2STD���1F�_��7QOF0o��5z%�2RC��6RC˰�86�"Q�bG�u 50�gMA�a_�q���QQآ�\B~�%eDIR�bGIvbqI�gaqG㓣HM��1C:�R� ���BF,SDN�Ҏq0?��MGTw1�`n�QL ��SMEf����M�U] !XYZU���AS�3T>���TRL_teKX��NU��!U-@kp+e�p�OL*fARE��S�I�B��ERWI�DT�$UPP1_!P�f1POW�\E�(�R���dS7�U* FTv�AJN�EM �~[d(V2_D_V_h_ �_�S`�f3`�P�k�Q��a�U�] �OV�4 )��AN \C1C�RW_I��P��)�h��h�K�p3�#��X4 P+;�r��?�,#v���im�D�C��WA2�AOT x$MY�΃��Xq o�fs�sS�F���D��x�����M_DO���H�LC����R�P��q��CU?�M17l���`���u�>�Z���PNT�V�PL�PV��#��!�p����@� PaXl�1b�BT������vƲ�uNS�VA�q.S�D	0Qj���Li'5EMA��1B��ENY}� ��SU�ZdۄS�چM�C)0LHD����_���Y�UZ�I�I,�I:� #�G.dm��|��|� ,�|�g���H�����f�EK�PI)d��K�����V�Rβ�CFUN�CM�����BBEL8W�L��AVIBj �t�7�� �&)�O��0�TRd�B�A��S��p�r��bS;���A�_D�F.�L��  2L+ ��J��M��å���`VRl��@YGLIN���q�Da�ߠ�1��H�`MG�����EV񑊤T!Hd�4�k�A�A<�ߣ&A�EA{�=�F� ��4 RC�����`DV����`F���P���	��CRTP<���e 2Np��csGU���DNYp�f�bPK+SA�PK�a��5��ѻGJ�bZ�DT�2��8��^�D C�%�W�s�c!$��� ځ�t%�j#��K@9f������%�����3C��f�SW"��EAh���B>�t���BACC�ADJ?�Fp�|1�$F��IFQ�.�J�aAF]��ARGgE_Lt���MOk�o$FS�!DS�`G@i@z�u���TPr���`_SJ1�0�Є�Q{2����*bY����DIߡ)����J��p�P�AM�C/�M�1�FU�23s��_J5���҃�s�Ct�@�CY_ P LC1IG1h7��J��4Mp��2INO7��$���CsDEVICE��Q P2`�&o��V�S���Pfg3�BY�l$?�O�PCCsHND}G7� R H;�GRP*�E� �b/�@��Uh����hB�$ CsL�  S|�g@��b�FB���FEN���&��CsX"NqT� d2`DO
�PM�9f%^AK�HOTSWjDdrV_SELE�Au�%q�Cs~ �BU T2`~�<dNK_x��&��[SHA��Z�#�$��,�20��'��@V� ���DL��U 
摺��$��0!;�J$�2X���3Y{q��TO�:s	&��CsSL�AV�p W  ��(�N���Cq_AuR	PUNqX $�OCPC_��B weL'���SH�P�@Y 4�Po�*!��B "?&%?&R��CF�bZ� 0y�ip#>a�`9f�`��5�aFIL���"s��$ID���$ �A,��#Wy0�&NT�Vt�!V
R�$SK�IZcT�&1<2D�r6J��17 C06�SAF{ �G5_SyV�@�XCLU�Q���2�D_ONL�,�m3Y#=ROT��HI_VA�QPPLY_WAR�31H�P�'�3_Mq��;$:�Y_A.��4=M��IOC_�1�6�CRC1�r�4%3O�됞5LS��$DUMMY47'B A��$} ��y &3 ���6|q���cE��HC,����UM��Dధ�ػa���AFsPCP�#�DTH��pEavP��NTQ���E,��B:��s�|"����$TRY���0�Qs�j#�0�� [  ���ART_����� �NOC� �\�MASTE�RoԁFYT�!�r!]� D��FP_BAΫ ��S!$�ђU_^0�\H�S����0��7  ^�h�cs��If�$!�2]8WSG�� ?_ � �a�`IGN@�'2a���p���lqh.b%fAN�N�jGMc��a�LATCH��`�0rj��g�d�R��bD�AY�f�>"r!`� <�q} �#BB�)$��#+C3'H'A��QEF� I=0 ga @A�ObIT�"?	$TOTA�*D��A*D	}�EM��NIb��mr�j��nqA�!�t�`���!A�D*�tr+C5r�EFF_AXI��%c&P�AՃO�p����N�_R��r!d��P�p��Â�E�i���u�PcC�IMqIy��q+�4�Ap��qr!e 0�aJ���yJ��1Z�A ���U�@po��CTRL_�CA� f)rT�RAN���IDLE_PWѰ5�F�I�R0V*�V_E��PeN�IAG0Qr!gw #1$�@| �TKЗ@����0��Pp��R��ݰAsVE�`����W2�$����9b�u�P�d���qOH�b�P�P2��IRR�	$gBRK��vAB��	A��
���R���  ఐ�*����Pf���S@��RQDW�MS�P��AXe� ��LIFECAL��.�L10�N2����;�ja0���C��icC�P�RMOTN��Y�� :aFLA�CjaO�V�aH�HE7a��SUPPO.P���a]�aL= ��ej�_X_2*ʥYӪZӪWӪm�`�>�䣍�_2XZ�6�Y2.�CO���PS�A��N��jap ��|��P�:RI��o#�h `�aACH�fSl����ev3m�L}A��SUFFIҠ� %���t�r+C�63A�RMSW��i� 8��KEYIM[AGMCTM�S�s��"���9a:ROC�VIE<�$qj ��BGL�$j`�#?ɀ�P��P�@p#k ���0EN���sm�IQN'��B��Mq�BK��JB�q�q�%ORI_CT�����:a� ���COF��t�EBU����Pq��	q��q����q����OF:��Hbl ��BƃOTh�5�8ң�"0P7_GA�TSCX��N��NI_4�j�R� h�զ0��I`ICr��O��ճ$�S�ē�M@������[�����A1�J`PqiqA��9�m_L $n�Do�eIo�T�`�$SKG�x�$�I�FBK_�W0DO��RK��@��AW_i�E@p�嫢˖@pz�SL���UPcCE�B䤯�LE�p�_��UF����I�T_�p��Ї������0#��>�1_�r;�]2A�1_I7�2Y�
�qB�n�rT�3T���BUF��՗�~֗�p�B�G�o�� U�<y�ղ4 �!@8�p)r}�IR�c��9�o����UP%an<P|m�܄q � ��T^�4�F�5LSP_���K�5���s4�1Ë3E8�!dc4�ARR��.�~�T���T�%`_�RD��5���SND�]�T���VSYP`D�Z��2l\���PmD��n-����Po���� pk���r�R���c+`��~����Pq �`�`���s�p$HOST0!�Pp�	p��4 ��p�EMAI�LXP��R��BFA�ULurtL�}�"�C#OU� :`;QT r!?u< $��%SlЦ�ITmC��!���DEVICE_9N�16�SUB��C�PC�$u��ek!SAVr%4"�M��1F���'�0.5�Py$%ORD=�Q��X%�A�(�OTTp�l�s��@L0���*1R�'AX�spb�0X��O3�#_G2��
PYN_��%pv��d;FDpp=D����쁠F�IF9`$U��POP�ED&�@EC�`�wMR�0	GH!7q&c�0iq�E_aNFO�x (�PSVv�.t���Iy�rP`wTy�p!��1��#C_RG��IK9bB&bD]�Rp4��1}��1DSP$��2PC`KIcyE�E��1�@U4G��&�CM�IPV��3p�l�VDCTHL�y�GE�pTJ�fWCHS�39CBSI�[���V�`ZI�sTly��tNV�@_G!�TL�TF��F2�5�d09CF�1:aSC;˕�CM��GFBCM�P�S�0ET��z6�FU��DU da��#�WbCDMI�@� ��� �EOz`}{�s!aI�@�Qe I��!�MS���Z��Pʔ�4�Q) A�|�� "�����4$Zx{��NIO_U<dd�{ePàwiCN���{`l�l�iGROU`�W�r���TMN}k  u�e u�e p||�i~cHR�B��bw��0CYC{�zsbw~c�/⡛zDET _D��v�ROS��q.fDAYav����vTOTz��w�tO�4��v�E�&�AL&�0ALa��}�2�!C��!ːBs�i��Q�RP�%�~~ ,@R8�%8�G�!LR�1}A0�0R AU5T�2�$�������˓$P�`��C"�@��O�5�A1��|� H��H *��LX��^`��VG�P ��.���.��.��.�P!�.�.�-�7)�8)��9)�2�+�5�1B�1�O�1\�1i�1v�1���1��1��2��2T5�B�2O�2\�2i�U2v�2��2��2���3��35�3B�O�3�\�3i�3v�3��3ʐ�3��4���@�E_XT_SEB�Q2���LTЬ�a0w�:e��0FDR;��T VEL�#?0	p��I⾲��LIFA�; +OVM�ܴ�A�TROV�DT} �MX��帳MO�0�IA� N	D"�ڲ
Nȋ0?0}�G'1ɱ�~<1ݱ�6� RQ�RI^�M�ܲGEAR�IO�ٵKԲڴNF���E�FF��P�0qܲZ�_MCMZ`����FEATUR�R�xy���J!? ?�F��? �?@� �	E��(��u4!U�����TP
q$V�ARIk�g�4#ET�UP2_ � ��3#TD�@��2$T��`8ю׈�44"BACK2� T�4"�4E)�:%�PB�"їIFI`�T��P�T�"@�LU��}�� вqBGLVܽC URS�TY�f$�2$P* �EMP���"$\�S�?�xh�J��� �#VR�TX��0x$SHO�]�L�$ASS��@�CU�@��BG_�������O���\����i�FORCn�pl�Kd��FU�	12�2�2j���@�"� |^�NAV�Ya�\����аS��N$VISIl��s2SC�$SEF�Ԩ�V Oa�$�\�а�p\�$l�I���f�FMR2���F ���P ur��� ����������P�����Բ_����?LIMIT_
��T�C_LMyƞϰ�D�GCLFY��DY&�LD8�|�5��s�P��B0��{�d�'	? T�FS� |�� PS0�3?0�$EX_1P0SP�q3<5<s�G!Q��� �^�6�RSW[%ONTP
ÏEBUG��ٵGiR�`a@UuSBK�a�O1��  P�O ���P{�M�n�O
t`SMo�E��"�@�s`_E ǎ 0� �TE�RM%�%i�OR�I�1 �%CaSMRpOm� �*AS)ْE&5�UP�p ��� -?�sbQ�\�##� �r�G�*� ELTO�A�p�0<PFI$c�1Ї�P|:$�$�$UFR��$���!� �UB OT7<PT�a��3wNST�0PAT�q=14PTHJ���P�E�P�3[p�!ART�c �%� c +2�"REyLu:�qSHFT�B(�!91g8_��R�P�SJR& ] $l'�0�b �����c�q�0I�0_�U�b �`PAYLyO�@vqDYN_��IЃB91.�Å�@ERV4�AR�8X�7S��u2����_Eߡ��RC�H�ÅASYMFL3TRÅ�!WJ�'X��T�EX�c1�IR��QU��DS�Ag5� SF}5P�@PC@Q�6ORS�ML��g�GR����	�@��80� uq��Hm��T� �?1�֧��P�OC�!�q�$OP�������б��dbRE�PR`�#�q��a93eB��R75�U�X1��e$�PWR���o�7@R�_|S\4^�t�#UD�Xӟ3SVSQQ�" ��|�$H��!^R`ADDR��H��G;2ka`aYaTi�R�y�m� Hp�SSCy���eߣ�eO��e�\�SE�|�QRP�OL � � \����bÅ�b�Z�S`UCLLV6tv�_1��V6j�a��HSCD���� $H�tP_"�p_�o�MrP?�>��LDT�HTT�P_��Hm� (���OBJ�pYb��$��LE*3�`�q�� � h�+qAKB_O�T��rSEP̒�,�KR�`�WHIT����tP��P�r��`X��P�ןPSS���'�JQUERY_�FLA�!+sWEBwSOC}��HW����!m��`�@IN'CPUP^�O���q�4����d���d��\����IHMI_ED~W T � x �H��r�$^�FAVh: ���N��RE�� @��@p`E}r��RQ�Lu��@DFY�U32$DUMKMY��H����!�IOLN�Ҟ 8�p�R��O�SLR$INPUT_��$�P��P��#�a�wSLAt �l�������vC��vBT�{IObpF_AS����$L�Щw���1�UR �0�!5�r�A�{�@H>���<���MQ�UOP�� `�Z���2�,�2�3����PP�3�Pz���3�������IP_MEܐ�ၢ X�IPx``Pݢ_NETPe�^{R������Q�DSP��{p���B�GP�`a�MaA"�3 l"�3TAB�pASPTI���E�� lf��0PSe�BU ID� �Aq���P��0�a4���+0���F�y�Z���Nٸ ڵ��IRCA_CN�� � ��y6��CY�`EA$��@w� �x��38�W�RS0x�A���ADAY_���NTVA1夰|�p��W5��|�SCA@�|�CL�� ���t�"����X2���N_�PC�����j�=���� �S,ђ���r뀌�fpp� � C3�Q�3���"���8c֤rc�LAB+1��\ ��UNIH�u�= ITYs�5�deԂ�Ro {���q�9�R�_URL@��$A��`��A^�n g�T��qT_UW�ABKsY_���2DIS\������J��ӡ�ؠ!$0�EyᓀRr�Q�"I A���[�JEqf�FL%����|��
�UJR��� ��pF-�7K��'��!���J7��O�B$J8��7Zo�����7����8���A7PHIt�Q�� �DJ7JY�+�*�_KE��  ��K΀LM� 7� <��XR������WATCH_V�A��!@�ѠvFIE�L�Vcy�U��խ� > !1V*@Ƶ�C�T������ LG~���� %�?LG_SIZ't�`� ��FDI ���  ��S�� ��� �. � ��A{:� _0_CM3�,�
�F�A�
��r�T(���2	�/ /��/. ;I .E�/ G9��RSx�H0  )ZcIPI��0�LN��j+R�f��DE��E�����js�EPL���DAU�EA`rp΀hT"	 GHiR����BOO�a��� C�ѠIT0W�G$��RE;�^(�SCR�s�DIr�S� �`RGI�� �p�,����T�"��	S�s�W�$����JGM�'MNCHL���FNK��&K7���9UF'8�0'8F�WD'8HL^9STP':V'8��'8N '8�RS�9H�@C;�C�Tt3�B�Rp�'�9U iq;4�'��%��$�.2G9SET?p�y:��%t3�4'�)9EX.�TUI5I^ � �^�r�C�#�C0��'$S���	��{%��@z!NO�FANA�uQ��AI��t���eDCSm��c-S�c*-RO3XO?WS�]RrJXSVX�(IGN ���)1��;�6TDEl;a�4LL5!���Ԡ���ñT1�$�؜��_�t3A
�������s���ᡭ��S1%e2%e3�%a,�bB.PԠ� ��{"`T��]%�����RqU�?p\&��fST�[�R Y���@�` _�$E�fC�k ��hp�f�f��Gc�Ԡ� L��*�� ?� � �c�p�h�rpEt���"^z#_ �\�ˀ�����{ ss�MC��� ���CL�DP[�C�TRQLaI��E�y�tFL,��r���s��D���w��LD�u�t�uORG�K��1�r��ERV ��(���(�Ƃ �s��� �耳t�5�tL�uv PT�p��	������RCLMC���(�:���4��1�M���h��b�$DEBUGMAS-�(f�W��U�$TP���E���N�FRQ~��� � ���HRS_RU���=q.�A<��5FRE�QP!$�  OVER{�)��_f���P01EFI��%�"q/���¡4�U��� \;�h���$U�e`,�?_���P)S$`f�	s�C ���U�����U� �?�( 	ơMISCΘ� d�eaRQ�d�	�TB� �� 1\��Ai�AXC�P�|l���EXCES�Ҥ�Q?�M:��Ѽ���P�C�_�?�SCf` O� H)�`�_Z�@Z�O�񫃯��=�K��a�ߒ�� �B_��FLICtBh QoUIRE�3MOO��O_�ǖ-�ML?pM�տ mpV!����t=����`MND��x�����!���۳D|��INAUT�!��RSM�����PN�{���3����ȲPS�TL��� 4��L�OChfRI��heEX]�ANG	R	�M��ODA8��L��ҧ�~�MF��5����i>r�@Hu�����S�UPDu;�FX^�I�GGZ! � � _�>s�!�>s�6>t�� ���bٵ` ص`/��0OC��W��TI������� MN��� tV��MD��I!)��3P�ԯ���Hq����GDIA��a�W�!P��a�A��D#)2��ODO�����4 $HW�N�B��N�TIN�aN �#pdI�ǖ�
���`-Lk SK�d������1�_Oq��!srI9 }pT�z�&�qFl���WAI�`O�t�KEA������>���V�aL1 I � �2��Mp�L$ae�j ��CA�LL_��ϑOR�T�v ��� ĠCU V���y²��� ��T`��^���R_NA�ЈEu��/��U�� OC
TR0`�p`�WMpIA�#��h��k"4APRbS�� M�P����ȏ $ F���3!�G ǖ��!_ꀽ�� �V`pc���ɒ����P��� �P�KE�2��$-�$B�� ND2x��r�2_TXGt�XTRA3S
<��qM���ې�P��`Yhf���s� SBp��eSWCSN��M<����PULS�S�NSr�J����JOIN���p��тr�?r��p`�т��?r��TA&��'�'�'%E�SF��RJ~�#6ePL$ ư��:e�¢DIR�OB�����LOAݢ�H¢�$��'F��e��&�#;�RR2C���h 6�!_PA����dE�Ib���G�!Q�'28<� �opRIN�@ 4<;$R0SW0��M3�<�ABC��D_Jp� V�	���_J3x6
r21SP��O@	�	Pr4�=3�=j�p	���5J<��5I��O��QI22��CSKP �zD���DJ�A(��QL8EE8E.Gf�_cAZ���1jAEL�Q<�2��OCMPtË��葱RT ��C�%1��G �%�`1ͷHY��LZ�DSMGRS�T��(�JGepSCyL��a�SPH_bP�(�	U��	�E�R�TERY03�(PA_L�`Y����P�c(��HTDI�A�B23Uf	BDF�jPLWoX�VEL�qINSrB�ApB��T32_���T�W�W�UY4Ѓ�0E�CH4r<�TSA_(Y1�PGdpT>P��`OFϱ��`��M�d`�U*`�MACC��M�W9 �@�T%��Epв�e�`e�p ��_ap_/� �me�bPU���d�"1ђi`V4 DH������ 0 $V 
0��S�@[��@~�Y��O��Y�N�RX��H �$BE`G�(Q_C`E�QC�3u�<�D�IRC_����T葻�$PS���rL�/su�s� VvF!0Vv�5y�wKs"�w3zr��_1b'����y��5q_MG�X�DD�qIRY�FW��ⵂ�Ks6r�D=E9�PPAB)�s^��SPEE�r[�j�IM.Ar���6qFbUS8�["��P��CTR��Y)�py� ��YNB� ȇ�0�YɁM�p���pO8�P�q��INC�n��8��i��31j�ENCY!e�	�rq6rg�op
C�O Izr_����C�NT�S�UNT231_mRr��LO~Pr��E.QD����PGd���a�Fe��Cx`t�7 �I��m �qĂ2CP�ERCH  HcO��.R �t��GѰ� 1DGѐG�B����W �3	Azrl�L���3��7�u�������ƖTRK,U�AY�#f���ۡ zr�ߣo��FA#�dpGMOM�%���Aj�j�T7��'���s~��� DU20�rS_BCKLSH_Czr m��떨�҂u�?������0ECLALM�q��� ȵCHK�
@���GLRTY K��_���$d!����'_UM��C%��q��A3Á�LMT�0_ALn��CL���W�EQ� r�d�P�gum�gx�0��0�w���P�PC�P��H��MO��CMpE`C`�CN_)2�N��3Sa@�V ����U�(Q��zrV���C� #�SHգ)2� G�$CcX��%{q�)�@f�PA"��_P!��_M@Ub�) 
A����J	b��\!xPO�G׍TORQU ���5ޓ��G������G�i�_W4�ۤ�A'���c���c��I��I
��I�cF> z��2��,�1	�VC5p0���T���1�����J�RK�H�;���DB��@M���MC�0D9L�a��GRV���0�c���ch�H_3e�����COS���@��LNJ�������@����@����#
��c�Z����h�MY��a�������	THET0��NK23�c��c���CB�CB�cC0AS�!�����c���SB�c�GTSy!��C�1��G����G8 $DU�򰏧].2�Ul�UQBL�_P�H��CE!AKħINX�`�A����3e����LPH������S�# # �/H#2*O�`EV�V��`,V*UV#+V1+V?+VM+V[+Vi)H�&2P-��%8#+H1+H?+UHM+H[+Hi)O��O�O�9.O*O�#+O1+O?+OM+O
[+OOF��-I�2D�SPBALA�NCE_q]C`G�p�SPea�B|�B PFULC�H`�B�G�BPrj1�'��UTO_��T13T2�I1r2NԱ�r ��T!a&��@��r,s�0�T��O�`Nqx�I�NSEG�rϑREqV6Vϐa�DIFǕf�i1�|W�b1��@COBrQ����B�2q����߱p�LCHWA�R[���AB��D�$MECH�q �,�Q�AX�P��f8��b�@� 
bf��*qW�ROB �CR�t�Je����C(q_���T � x $WEIGH�FG�$��c�I�櫐IF���LAG�ւ��SւaPւBI�L�eOD�Ґ�bS�TBp�bPaQ���`4Ppu�jas`�w`
;�x(rׁ��  2�ݔ^�fDEBU�cL�pz�b\MMY9ju�`PN��KtG�$D��q'�$5p�� �	��DO_:apAra� <�`v��@�ׁ�B�b�`N�q��x_��׀�bO�Ű �� %")�T^�f�9�TsQ-t�mpTICK�c�PTE1up%�sd��N ��@�s �R��ׁ�R���R$�|pPROMP��E� $I�RI�Ձ��_����MCAIm���x�_�`Cv�P��R|�7COD
sFU݀�fID_����_PY�e@�G_SUFF�� ��ć��D�O�VP��`�GR �c�R��9���R��R��r���|tpֆ`Hn�P_FI	q9n�7ORD�a y`=r�36��o�Ձup$wZDT��	E �a�u�4 *�QL�_NA�q�Ȓ�DEF_IؘȒ>�� $��b��d��$��>�IS�JДq���DW�$��]�;t4ф���bD�@f���
sD�F�Og@�rLOCKE����*�<�Y����UM��Ȓ����� ���e������� .���fY�Y���P�� �Ȓ���`�����pP�PG��pS��mp�W٨صϣdaTE|ñ�t�( �a�LOMB_��0�bVIS ITY�bA�O�cA_FcRI�C5åPSIS��7��1R�^��^�3#s�bW:�WF�x�<�rL�_���EAS�c���4ģП�~�_�4�\�5\�6�cORM_ULA_I����wTHR�b��G����w`� 3|8CuCOEFF_O�qMP`�$�q!G�ѢcS�`\r#CA�@ass$�ác�`�aGR� � � $Ϡ$R�rX�pTM§��ϥ�rXף�ܦsERpPT��ܷ�h��  �BLLt���S�_SV��F�#���h��U 5�h��� ��SETUS�MEAn�׀���`��ao�s`� � ��;` :pг� b�᧡��͒���á	������$���D����n������PΒ�REC���� ��pSK_h@���� P�a1_USERQ�RL�PQL�QVEL��L�Pt�h�r�QI���@�MT�q�CFGB��  ���PO�RNORaEq`�p���SIra1ߨ�v�RUX�����YQͲDE0 _$KEY_(s*P�$JOGT`S�V7Ua����SAW�R=�����T���GI�@e`OPWO}R� �,ip�SYSBU� ��S�OPu8���T�
U�PPϠ��PA`O���R��OP��U�Q��Q��$�� IMAG��*P�� ��IM�IN�����RGOVR!D� �P��P� �@G`b����I�RL͠�BT���PMC_QE���9qN�0Mx�Dq=r1Br��(SL��@C�� � $OVSL!����,�"��2�REPq�_(� ?�)�?����=r#C8`ʐ"#!�)/_ZER�����w$G�� ��|��B�� @ ?#�eORI��"`
�}&���)�!�!��PL����  $�FREE��E\?���PC���t� h �d���w~��PWR_WS����EN5	1REM88%5	1HWH��3�?41сQE'!C�� qH�a�P�`ATU1nSqC_TDXu6B�Ђ6k1��}�CqW3��C�� D�q� �� �0T�t�d�"�RXE|0���2�2�4r#1�y �`{0UP��o��M�PXb��6�;t3��2� G���8�SUBj1e;�j1��#JMPWAITX@��ELO>F�qS&RCVFx�	��R��ARE�@FWQ�qC�& RL�R	��GIG�NR_PL�#DB�TB�`PQ��QBWȦ��D��U�p�EIG��H�I�STNLNl�F$RRT[NO��yNH�%PEED@>�HADOW�`�S��ERVE�vT��8TA�SPDB�� L�``㑢P��TCUN�`EK�P'AR�0�.#LY���@1cbP_H_PKT�$��?RETRIE�#�����Uk�FI�"� �y`�P*d 2꾫�DBGLV�CL�OGSIZ��K%T�AU>�gdDaS)PS_Tc"��M�C!�&�`vmR�c���B�HECKP��L�9P��Q� 0{ h�`qAL� ��NPAⶠT�R't��PIP4�#�P��"ARZb���0d�+�\0O��B�ATT�p@+�Zf�`0�r��Es�SUXd :"p8�� ����� $��9ITCH}B��W�O�!�#�qLL�B�Q�� $�BA)�D����BAAM� U���v�!�p#J5 ���r6��q_KNOW�c�,�U��AD�x�ЭPD�O�<�PAYLOA��`�Z�_�1c�xc��Z3L;�1� L_� !{����q���=��F��C�����⚄I�I��R ���~��0��B���3_J%!�_J��g�=�0TAND��`?������!��PL�p?AL_ �p�P�A��Bk�C��D:_�E���J3T�h��� T� PDCK�dP�4��_ALPHx���BEu�2�x�Ɗ����Qb �� �b�Y�D_1j`�2��D��AR54�>�(�L�7��0RTI�A4f�5f�6��MOM��r����������B�@ADr����\����PUB�R�� ��㥌�QAC�h�%���P��"�i�aP����R�q?��� e$PI!=Q�X�e�P[�!�[�Ig�Iu�I��#����8A��CA�0O��V# %ZSHIG�sZS�E�T���T �E�@�@��3���A�<�A�ESAMP�0�a�j���pÚE�pE� O����M��8@��ƟP)���7�MRO��1m�Kd����KIN��d�S��!��ĚB��G��G�g�GAM�M��S~10rX"ET��"F[ �D���
�$k�IBRA;RI,~AHI��_�0$����Eސ��A�����LW��$���H�����1Pj�C�EC�HK6� ����I_R�<p��>��c���ű璣��Ԧ��h� ��$�� 1���I� RCH_�DV���aS+�LE@��X�!=����>P�MSWFL�D�S;CR-H100�c`��3nb�����r���x���P��PI3AJ�METHO:#���EV��AX�#�0X]P���;RERI��o�3���R�P5�	�$0FH��p���P��B�]	L�p�rOOP�����APPK�[Fb�`���&��RT-g�OS��P�e���2L$�c 1��Z$� ��RA��`MG�!2�SV�>��Pp`CURx�LGRO`P�1c`SA�qONnbjCNO$0C�! B�j ���k�}��������2���(7�DO�QA �ҙa�Ũ�����q��q3�h'd%"#�� ^VP�$$C� S(p���� ��'pf'p � ��SIp�&� Y5��ܐVM_WRK� 2 �%� 0  �#5�!�/8�/)= )<	L0==`?�'p� �N?�?r6�5 <<�=�?K1�?�?OD�� BS�;� 1��)� < �?UOgOyO�O�O�O�O �O�O�O	__-_?_Q_ c_u_�_�_�_�_�_�_ �_oo)o;oMo_oqo �o�o�o�o�o�o�o %7I[m� �������!��3�E�W�i� Bh�c�LMT� l�d9C��~��IN�����}�P�RE_EXE��ր��_UP�ʁ1J�!� DV� ST {�'%?�*�J0�Q�HIOCSNV�ȕ�Pl��USʅ5Gi�_q� �1�+P $�0�`v1ϝ�<̟� ?�Z� �����%�7�I�[� m��������ǯٯ� ���!�3�E�W�i�{� ������ÿտ���� �/�A�S�e�wωϛ� �Ͽ���������+� =�O�a�s߅ߗߩ߻� ��������'�9�K� ]�o��������� �����#�5�G�Y�k� }��������������� 1CUgy� ������	 -?Qcu��� ����//)/;/ M/_/q/�/�/�/�/�/ �/�/??%?7?I?[? m??�?�?�?�?�?�? �?O!O3OEOWOiO{O��O�O�O�O�M~�LA�RMRECOV �텰�����LM�DG �Z�~-R_IF �����d  RVO-�002 Teac�h pendan�t E-stop� cation �error ,70200408Z� �_�[pP�_�_�_o"o~0j, 
 0o�Yo��8ROS2 ~vjLINE 0va�AUTO ABO�RTEDvhJOIaN���o�o�e$ra#  �`�o�m�e�o��\CIuP20 L�BL[1] ex�ists in �line 1:  0 tew���o�;e	QWAYS_ON_DO�����NGTOL  �� 	 A  � ��~�PPIN�FO 7[ �VJ�\�n�����  Cb����R��ُÏ �����3��W�A�g����@�����˟ݟ ���%�7�I�[�m�������)�LICATION ?�u��D`�LR Hand�HpgToolvc �
V9.40P�/55���
8�834�b�240347�2����|���7DF5��vcNone���FRL�� �ub��*�_ACTI#VE�t£�s���`�MODɰ;e�yP�_CHGAPON���q�OUPLvp1	_Y� <��@�R�d϶�CUREoQ 1
_[  �zn�n�	����Ơ ��S�ϳ�����������g�1�R�n¤ԥ\�H��u?�r�HTTHSKY��R��\R� d����F� ��$�6� H�Z�l�~����� ������� �2�D�V� h�z�������
���� ��.@Rdv ������ *<N`r�� �/���//&/ 8/J/\/n/�/�/�/�/ �/�/�/
??"?4?F? X?j?|?�?�?�?�?�? �?OOO0OBOTOfO xO�O�O�O�O�O�O_ __,_>_P_b_t_�_ �_�_�_�_�_�_oo (o:oLo^opo�o�o�oL�o��TO�p˿���DO_CLEAN�Ͻ�CsNM  �{ nϑ�����t�DSPDR3YRJ��HI�m}@~E�W�i�{����� ��ÏՏ�������MAX��*t�a�aǂ;�X*t:�7�:���PLUGG*�+w7�۵WPRC�pBkpo{4�&���O����/SEGF�K�� ��k}E�W�i�{���ş��LAP"�5��� ����)�;�M�_��q�����������TO�TAL]�3Ɵ���U�SENU"�/� �xϽb��RGDI_SPMMC��љC	�M�@@�/�O� �B��+�_STRING 1���
�M��S���
��_ITE;M1��  n���� ���������"�4�F� X�j�|ߎߠ߲�����������I/O SIGNAL���Tryout� Mode��I�npL�Simul�ated��Ou�t^�OVER�R� = 100���In cyc�lR��Prog� Aborh��~H�Status���	Heartbe�at��MH F�aul����Aler�����1�C�U��g�y�������  &s��&q�ϲ� $ 6HZl~��� ���� 2D��WOR���|�� V������/ "/4/F/X/j/|/�/�/�/�/�/�/�.PO ���� 0�	?C?U?g? y?�?�?�?�?�?�?�? 	OO-O?OQOcOuO�O�O2DEV#>�@7? �O�O�O_!_3_E_W_ i_{_�_�_�_�_�_�_��_oo/oAoPALT��ha�Bo�o�o �o�o�o�o�o 2 DVhz�����VoGRI@���� �o�4�F�X�j�|��� ����ď֏������0�B�T�f�x���R ����$���؟����  �2�D�V�h�z����� ��¯ԯ���
����PREGlnU�ȟ.� |�������Ŀֿ��� ��0�B�T�f�xϊ��Ϯ���"��$AR�G_|D ?	�������  	$�"�	[�]���"�8���SBN_CONFIG���V��U�o�P�CII�_SAVE  �"�x�k���TCEL�LSETUP ��%  OME�_IO"�"�%M�OV_H������R�EP��!���UTOoBACK����r�FRA:\B� ,�B�x��'`��B�u��� �����24/03/05� 00:23:2�8B���26 05?:36:02����52:1��9�B��hꈄA�h�z�����X����B��!`�_D�_\D�02\W�SLOG.DW� �2D��`�CRXL.Dkl�������V� $6 HZ�~������� �  ��A�TBCKCTL.�TMP CFG_�RPT��PEAK���_OUTPUT�.V�G/Y/k/��X��m�u�>�INI�k`��h�|�A�MESSAG�Ж!x��>�+ODE_D�ЋֈhՉ$�"O�@�/>�PwAUS40 !��� , 	��9��8?F7,		 0?j?T?�?x?�?�?�? �?�?�?OOBO,ONO�xM40TSK  �=u�/�A�UPD�T� �'d�@�&XWZD_ENB�$d��FSTA�%��E���XISV�UNT� 2�Fu�w�� �	 �/ �rW. ������� �� ��ΦB�PP����*��u���k_�_��^PQOK  �k�Wֿb i�� �#u ��ѓ_�_�_�_*o-VM[ET��2>Y�w��POQA8�y@���PA 3�?h�Ա@?�A&�cm>��=�v�_>�7�<���+>
P�<���3mSCRDn  1�W�' ���u�o�o �o#5Gn�B�9� �o������S ���A�S�e�w���؛�����$D�GR`7P�@�/҃��NA����	D�φ_E�D� 1�i� 
� �%- ED�T-����P�t���Dw���-D�C�B�9�A7���<��wp�ܕ2���ß@��D���@y���ҟh���ޓ3�� !���E�W�گE�����4�¯ޓ4}�U�ʿy�2X����X�j� ώ�ޓ5I����W�r�@��$�6���Z�ޓ6� ��bߩ�W�>ߩ������&�ޓ7��Q�.�u� W�
�u����d���ޓ!8�ﹿ��ݿ�X���@A����0���ޓ9y�������X���T�0f�����ޑCR�� ��R�l�0��TҀ�NO_DE�Lޏ��GE_UN�USE܏�IGALLOW 1��}P(*SY�STEM*z�	�$SERV_GRp�z��0REG��$�z��NUMx���PMU=>z�LAYI`z��PMPAL|� %CYC10�1. .W#ULS�U/�3"1�L�m/�$BOXORI��CUR_� ��PMCNV&� 10G.� T4D�LI�@�/�	*P�ROGRA�PG_MI.I?[0�AL)5h?R5[0B��?�$FLUI_RESU7'�?���?�4MR�O
�SET��DATA�-O�$DPM_'SCH��� R �O�O�O�O�O�O�O_ _+_=_O_a_s_�_�_ �_�_�_�_�_oo'o�9oKo�	ҀLAL_?OUT �����WD_ABOR�8 aс�`ITR_�RTN  z���j�`NONSTO���d �hCCF�S_UTIL ��ʇCC_AU�XAXIS 3"{ h{ohz���čCE_RIA3_I^�e�pn�pFCFG �"}��$��q_L�IM�2)��Xp� 	��B\��z���
  .m�z��Zz����'� ����Y��`@��,"�������u�J�z�
3����1���`<�#�L�r��PA�0�GP 1F|�s�����͟ߟ񟰖CZaC��C7�J��]�p�����W C���+��+�U���+�����U�+����+��+�e��;�� Ck#��+��+��+��+��J+��+��+�J��+���+��� D�W D������m�� �޶?�5r�HAINFAILKDO�f)w��E�ONFI@�o��G�_P� 1F{ )Fu(�:�L�^�p����������KPAU�S�!1Fu�s  G"���Fuܿ� �*� P�6�tφ�lϪϐϺ� ��������:߰��c�A=�u6qM�`NFoO 1���� �1�;����?�?���>N�c=l>(�M��3҈��t��@��A�9�$�`��@���ڴ� ����CD2jD4��
Ca�������v����p�O�q ��x#�L_LECT_�r!���6qM�EN)0�eiܬ�#�NDER�#��-w1234567890�� Y��������ЅzByo  )�*���� o��H�Z���~����� ��������C 2 �Vhz���� ��
c.@RЫv���$Z� �g��IO &�阅���f-/?/Q/lc/�TR��2'�Ĳ�)
�q.�(�
-�*�n�_MOR'A3)F}���$51� $9<?*?`?N?�?r;�"T��1*F},�?������3��K�4��6q%P��,Z����-O ?OQOɏuO�O�f`�%���@�܍O��� �sja  �!}1I�PDB��.��l�cpmid�bg�O)_!�;S:�ĐQp_n_9V  ��_�_}]܏_[_�_}]/��_!g�_Doo�^f3o�o�,ݑo�ud1:�o�o{��ADEF �-$�#)�ac��Qbuf.txt��o3\�o�0�/���>��|2"!Ry�MC220�K�dX�u�s321�}��t��u��Cz?���2�B�GGA��{A�:L�@$��A?"��B�������_CX�VB��JA���B�B�C���Q��EŚEM��Dfn6C���D��E�d���>L�͝�Xs�623�,D>�����U!c`2���P�c`5�C
��x����}���  D4��C�����  E%�q�F�� E��p��Q�F�P �E��fF3�H ��GM�8���?��>�33�~�C���Hn���A@F�B5�\�t2�@A�1���=x�<#��%�# �O #��-�QzRS�MOFST +xzH�V�P_T1as�4�-A ���M�ODE 5�= � 5���!���A;壞�����?���<�M>�y�^TwTEST�b2~���RT�6-���vC��A݀��	� Ӂh���r	�C��B�,�sC�@��w����:d��# ���Z���Z�r�\�ϡT�_�`PROG �%�:%D��̤ N�USERi�ѵKE�Y_TBL  ��5t����	
��� !"#$�%&'()*+,�-./��:;<=�>?@ABC�`G�HIJKLMNO�PQRSTUVW�XYZ[\]^_�`abcdefg�hijklmno�pqrstuvw�xyz{|}~��������������������������������������������������������������������������������͓���������������������������������耇����������������������[ё�LC�Kۼ�Ҵ۰STA�T!�ͣX|�_AL�M߸���_AUT/O_DO���vӿFDR 38{2�`�AX�q� �EUOSYS�T-325 Pa�yload er�ror is d�etected �792004017,70��0 ������D$JOGGI�NG��1��MF��AC1��=���B�	i�A?���`�@���Ә"W���ΨC�@q�C��<�{�w�;�� �B�P�� B���J�@� ��� Q�}������ C�W�H��1��CB���B�z�p�X�R���@��0 Cont�act forc�e exceed�s limit �1,��Y���� ���2G�'� �=�VO�	jM�A?��`���@���c��Z��C��C��$�>a���=g+�oB�̂��͈xqR��F��� �� ڠF@���G�����I�������8��a�s��������G�3�������@����A�>�`���@��xqf�����CD1�D4���=��77�E�B��*�‫�b����7� �R� �{�����p2� �� �o4FX�A
�5��{������8���J/���������@�+�|��1�&�CD22D4��n=&��"�ӣB�� B��ȸJ�你�����oj������6��X�zu�-�?�p?#/��?��?�c V������sr �A�{9"�@���!z&�� &D4��Pz9)��B=���/+ �pY���_���(�p.��ߘ��+MO?�fE70v ���/�?�?_�9���8t �0��0!���<��4>AvG|�C��WvO )����Ҙ���Q%@����!�$�SOeOwO���70��O�O�O`�O�O5/fo��V��=%f�0;_�2%�0�ZwB�G�B�I��T�-��U��Ę���,�pJ��ʧTr�_��_�_����Xz#h9;?M?_43g?��Kj��VA-�� NK1B߀��A����e�j?��§�� ���>c� ��]D9nC��߻B��d�v���C-��Ђ�M}-��o [;@����! @���O ?4&5�X{][m_?�����O&��8;S��r�w@j�����3?ܤ��^K����c�B��D���C���<�E�Ew�����A�9F_�/��/��/��;@/�����$�/��o�����
e	��p��͏ߏP������m <\7�G�5��(���:�@�¡�n�%���c�)��C����C�c�Ctv��סB��B�U�� >�:h�������CA�XV�h�ڟTK����t
��|��-�?���c�u�濙���3G���"�����{@��*¡Z����nc�YC���C��Cx|�:7�B�PYB»%'��58��� P�g����3�(y�W������{������1���Ϳ>߃� �<��B�e�@�-���yd@�S^ ������c�QQ�D�	YqC�zC�w���1��B�����VZ��
 P� P�c���ߔ�P�߸�Rr�t����_ocb�,������T<��X�=��:P� ��v�O� ���<�ӈ�8�C��G�C�B=����<\��Bw�ߊ�_�O�C���$�a�ڃ��a�o����&5R�� X{^ ���ϟ����︕�X>h�������|*@�P�����σ�?��C�I�C期�=Q[W���{Ҽ��@,��W�� ;;@L���� P� ��Α��L�^�p�"9����;�M�_�q������f	y{��b��!� u�7 ������˃�>��C�J/C�l�<��aX��B���Q Bn\���� 1	G���� P�AK��������1C�U�/	}�x��� �� v���*���?6O ��%n�39QY�B�.�Q�q*���G�Γ/ /0/�O����[/m/@/�/�/�/&O	���((� ys��U��̓�=�O ����R=3� wB
��B�ޱ��P�-�K?�� P�-N���vh?z?�O���s��������P_OOl�_9I���'l��_@G������<�C�H1��:�>^���Q=t� B�~2�8YԫO�bA���ً�@@�o��O�O�O�9��%_-_?_��oc_uPJOGG�INGMo�o>�G���g��0�� oY@Q!������ȃ׿'C��/bC�J=�}q7q<H�B7�uᇒ."����@@�@@�G���@ˑ�O5o�oYo����+{o�o�o��o�oF���?�S����3�� n�7 �����u�bC����3p�=c��5���B����g���O��J@@�@@�kh��G>P������.����p�#�5���Y���g�:�� pȊwд�����
�������TC��>�����<�Q�L���~�x[��@@��a"����(� �4���4;�M��_�Я�����Y�)�|ǔ. /k� �6 �<�����>~~���C��f��߆>�7�W�m�ߠB��`4�=���f��_��@@�@@�_�E�W�ȿ{�����;������0�����f�Y�D+ǔk���'r� ~�@WE���\?��C���C���C�߆=@�ڷ����B���Gr�HI
o���ӿN��{q�����r�ٿX��@p�?�?�3�4,70�2A8>�G�Y���]�P������#� {_@HbېR?������Ü�=&��;Ү�xRB�SLk��%� W� IIkfxw��� <G���&�8�p����\ �������u_&��X�?�C'q���� yH��ې��W=C O �s@�>?-�&w�>��l�B�gb� A��gw� L� FB@@�'�S��nqt�f7t���
Y� ] ������P���9����^��7��� `�@V��ې�_�7@uC��K�C椲<���n�;����B�h����U�T����9�[9�D�v�<�B�f?�I��� a-?�cu��9�Ȼ�i���� �8@IV�ې�_�7;AC��G�C�U?�
6�7!>�y�B� KGr�߶&7 >Hq���G6D	3�@@�@@�/AS j{��`?���F?Y��ף!�B�1h�Z����0=�?���� �9���A�SC�ն�C�;�=�����1<�nB�Gݜ��:O/��Ԥ@@n�R��@@��,�~�/�/�/� m �/�/�/pO#?5?�OY���cǒ hv����M+X?���~�d���J�IcC����C���=1��E�A;�X�Bw��C���rw�?+ !9�T,`��T�9�kaێ�?OOji o;OMO_O�_�O�O�o�@�D:��	4��L�>?���7�@������G2C��=�C��D=�a8�Wa<��B�C��G"��:�?��
���9�Sn�<禁�b�K_]_o_�/9� Λ_�_�_0�_�_�f�A[g2����A��������y}#¢n�YA�"��B���D;�C���=�B��q<��PB�A� �76��oo�惱����o��o��oX�,y�o��C��Ə�m"��p��A�����O��y`¢m��A�#�w*D�;`�p�<�������B����;�	�������9�_q1��2<�A����q�a"!����(%�7�I� W��[�m���🣏U&����4g2�
�A�f�����E�Yl�8�PB'��@�v��DK,�OC���=�Q��w�<ԅ�B���8�� "/��	�g����3���#u�(2����!W����͟�ߟP�����ɩ�G��A�e�����M�Ya.[�2�_�b�k�mDK+��C���>��,�ױ=��B����2?Kb�����*���9�5�#o"䯠ʯܯ���"W�� �-�?���c�u���)��e����VA�����&��*��G¡�BT��Y�C��*DJ���C�
�>�� $7�=ׄuBw��
�������0̳�S��6<�FU��2�D�V�(K#W��{ύϟ�������F�)�i��8A���t��*��*���г�a#ػ�DJ�CC�	��=Ď���<��ߋB��%�q=y�6
����0ܵ�	 s����*Ϝ߮��߳�W��������p�#�5�����t�g2�QP�A�7�3A��-L�м�Z�#ֶ�D?Ξ�C�M�>������=��{B���~! A�����)�Q�4����0���w������%W��;�M�_���������0���A���2�B�-�DDЖ�T�����D?ϵC�T��=	�W{���W{�W E�t2O��vd�0 ^��:Qn�Tfx�)&W�ț��0/���f/�銌��R8�AÐz��.��,�+¡��Ўa&ӵ#�D<�НCĸ�=)���"� B���gb= ��U���Z�0��0��9�0���������W��u'W���/&1�>/�?M/_/�? ��䧲�0�A�����9w�-�q� D?�ID�D��C�>��YA=Y5��B���G҅�.V�/����9? �Q*�$���[D�8?�$?6?(�(X�]D [?m?/�O�?��&_و������CA~�}��,�4�������(�BH��ѣv�LD���CQ�>O�a�wQ=���Bw�d�G�m�KwO ��)�t��8o�@����|O�O��q)�@F�O�O?Po__�o�9Y��GTA~y_]�,�TWPh[P�S_P�cW�D��C]�>7���a=�zMCw"��1/OK��? �����k���fA�c��_�_�_�j��*X�m/ o-o�O�co�?�������GR����Au�������i�QM��A��I��A�C�D��CSL�z<Ҩ17�0���B�����w7 ��W? �(��3J? �gO9����_��+X蒤 {�����F����0!$��C!�Awx���i���Z��A��BA������C�ECSR��<�ᗑ���{��� @�*��� ±X��-�$��n��ZB�_��
�����,X�T{ۏ�?op�#��5����x��rg�1���=���	�i|A?��`��@�������ΈC@q�C�?�<t ��X��Cj�X�>
�U��o�?Q�? �������k��OD�-X�qw;�M���п��x���D��+�ǣ��=�CӠv�נ�۠ߠ��ׯC@p��!s����*{�T�W� !u�"ѮW`��C��U��y����.������E��5 Pay�load err�or is de�tected 7�9200401,70&�8޿���j���J&Ľ�=ꮥPӠz7�颺�.�����5��r�A�2M����8G�@'��ϵ�q���� 
�E/�������8/��A�S����N���=W��Ӡ{נě�kδ�Y�ދ�oB�M1����? 	���<������9�C8A0���������`�����&�fǤ_�=�ǓӠ���風������F�A�unq�`��v��S���n�����$��8A1��Ż������P���CF�Ǥ�=�"@	i��נ�۠?̙����N5���B+����!D��`�� ��$�!4�����8C� �$C�R_FDR_CF�G 9?Q?Q���
UD1	:7W{�j�$�F&�%�s"HIST 3:��%#�    ^4_҂� �Q�P�_��_*q��_F$_dnq�`_�`_'�$�/�_7M/I?s"INDT_ENB�S�"�.�s"T1_DO%>Pt5r#�T2�?�7VAR �2;�'�P t�RE/d��?�|�?d��Z[%��s STOP�i?{2TRL_DEoLETE�6 [J�_SCREEN ��%t2kc�sc �!UL@MM�ENU 1<�I_  <xl%xo �O\��O_(_�b_*_ c_:_L_�_p_�_�_�_ �_�_o�_ oMo$o6o �oZolo�o�o�o�o �o�o7 FV h������� 3�
��i�@�R���v� ����現�Џ��� S�*�<�b���r���џ �����ޟ��O�&� 8���\�n�������ʯ �گ�9��"�o�F� X�~��������)�C�RE~ =�)�2X�T�  �x��� AA7A6?JS4125<@�C_MANUALPOn{2ZCD|!>�9��2e� ��"�Fn"d���d�?|(����dr�GRP �2?�9� B�����?g�� Ҟ���$DBCOb0RI�sEs6�G_ERRLOG @�K�!��g�yߋ� ~�NUMLIM#�1dt5
�PXW�ORK 1A�K�V������!�3�N=D�BTB_fA B�C��#��q���!D?B_AWAY�30�  GCP t2=s�׽ҋ�_AL��d��_�YO@sEt0�v6��6� 1C�� , 
��� �"�C�M�_Ma0�!���@�[�ONTIM6pG�t4�}����
����MOTN�END���REC�ORD 2I�K� �K�L�G�O� L���?Qcu }��7�� ��F�j�� ���_�W/{ 0/B/T/f/��/��/ /�/�/�/?w/,?�/ P?�/t?�?�?�??�? =?�?a?O(O:OLO�? pO�?iOO�O�O�O�O�]O_�O_H_�NDEXI_�_�__�_�_�_�_�NP_C�_$o6o@�_ZoEoSo�o�N8}� �o�o�oNoro'�o K]o��o���8���#��V�T?OLEREN`k�sB����L����CSS_CCSC/B 2J��z�� 4�L���Ώ���U�� (�:��^�p���Q�����L��������!� 3�E�W�i�{������� ïկ�����/�A� S�e�w���������ѿ �����+�=�O�a��sυϗϩϻ��� �ڟ���L���p�LL{�K���r�P�� CL�C�p��d�L�|� A�a�%pa��������� �? 	 A������B���?�  ���B������z��aL�B�L��g��m�P�ӏ��L������������L���(������:��5:� Ժv���ȧa��L�Ț� �ï����E=��0�U����&Nh;=���=���>B��RW�ȝ@��� <`+H;�?��<h��Z�����Ȝ��Ad���d�kA !Dh�Dzu���������W'�B(x�_��������K�Pؐ`�0�;C(  �� @��
�nU�i�oț k�Dȓ>m���C��a�� �[�YR���рXZ�ȗ��%/�/�I/n/�/�/ȗ�CHa�t��u�BB�?� D� ?[��/�/9/?Hu��!L�??��2[4�J9�=��w1<)�.��?!�F1�3 �݈3�7�9�?�? O�?@�?OO&OoO��� ~I0OBO�Oȕ�O�O `��I�/!_3_E_W_/ {_�_l_�_�_�_�_�_ 0��dЧ�0hw\ ���=uB��B�R@�w��?�;��q�{��A���gH��=8��=��o=�����Єo�o�oȞ�R���@RțD�@�J�@��@lx�@��@���@��o�B}�d֤�@��b�dN�N�d��Yҳ�d>���@�*�d,�@��@�GY�Tnq�aK�@��@j�d�8�@��d�Yҧ�b  ��@^�vq|�@��@��Y��Ш�rN��dN�@�R�d��Y���t��@E��@��d"�q�/�*Y�/�@�tt~J"q��d�g�Y����qFq�q��	wt��ts���ց�'t~[�@(�d�ۏY�u���q^q�a~��d����c��U��@�@��d7wr��P�N(��!�`w������v��1�t��*�g�����������$���C����QA�x A��� A�8 A����� A� �A�辐Ր� [A齐�`ΐ`�_����  H��F7230-0?003-01�*'� 9�K�]�o��������� ɯۯ����#�5�G���R0x13?1EEE70�-{� ������ÿտ���� �/�A�S�e�wωϛ���VR�����&� � TS120�-602-1c�//2B3Ab�2~��av�C2�159��/�06M�C�087�-901.�17�993]�o�035}�/�3����2���V߈� zߌ�>��v���O� �����G������� ���)�;�M�����H����u�
��P�
�� ���6�$Y�y� ]
�����&8J��ne	  V3�3��#~]��C4� *� ��� TT�*P��C~�C�� {�P�T�X�\�h+����~�Ä�L��A�r0>
�@��/%/7/�)nO=�((Q��Ui��!����$;Pz�ɕ��*�u0N	�=���=!!=06�_<CD<&��<�^;z��O�v�����B<]y{;�M~< ��s�^�O�mPA   x�/�+O@�  ?�;2Q����Ps0c�BH�V�X��0���=E�A�K�@�B��X�W�gz������A8��S�C�ܛAC����?jO�?�c	3>o�{�
�A���<`@@�$<`�2� Bf�C>�3�1C��0癙�2�4<��o?�PH�)S�B��4,1�1��2�0B��?5Bw����@����bi�A(�?��0r�D`oE»h O�?�OSC���@�T��b0�A(���0WoN �C0��!�� �§2	C:C\�2�`�B�?�0�Uo��?�����4��
m�$DC�SS_CLLB2� 2OoEf:0<H�=���"Qz��P�_�%=0 �n�P�_�?�ja�_"o�`�1R0 <@�"F�"�-@
 @A@A�agno`�o��o`�@�o�d�o�d�>L9P �2(V3B�?�@A���PD�P@���?�33�aC~Q�/�RV�@?yCa�9d?�0<a��VV� �1�AOE;� �u�AŴp8�u{t� �cu �����a�	� ��-�?�Q�c�u���� ����Ϗ�����)� ;�M�_�q��������� ˟ݟ���%�7�I� [�m��������ǯٯ j����!�3�E�W�� {�������ÿտ��� ��/�A�S�e�wω� ߭Ͽ���#�c��xTX+1aF< ����aư�����o�� g��ߝ�K��������=s?���_�����������C�&LDCKREC�M�a�1���)�JY���
sF��oIoJ 0���	��8 \nQ����� ��}���qC�D�� �������� ��/.//R/d/G/ �/q/�/Sew �/*?m/N?`?C?�?g? �?�?�?�?�?�?O�/ �/�/\O�/�/??�O �?�O�O�O_"__F_ )_j_|___�_�_5OGO �_�_}Oo�OBoTo7o xo[o�o�o�o�o�o�o �o,>�_�_F� 	o_-o��#�� �:��^�p�S���w� ��ʏM�q��� �Z�l���������Ɵ �����ߟ �2��V� ُ?�����!�3�E��� ��;��.��R�d�G� ��k����������ǯ ��*�<Ͽ�]�㯄�ǿ �Ϻϝ���������� %�J�-�n߀��϶� ��Kϡ�o��"�e�F� )�j�|�_������ �������-���T��� )��ߜ����������� ��,>!btW ����?��c�u��� �:}^pS�w ���� /�$/� 	�l/�%�/ 	/�/�/�/ ?2??V? 9?z?�?o?�?�?E/W/ �?
O�/+O�/ROdOGO �OkO�O�O�O�O�O�O _�O<_N_�?�?V_�_ Oo_=O�_�_3_o�_ %oJo-ono�oco�o�o �o�o]_�o�_"�_�o �_j|�o���� ����0�B�%�f� �oO��1CU�� �K�,�>�!�b�t�W� ��{���Ο����׏ ��:�L�Ϗm�󏔯ן ��ʯ��� ��$�� 5�Z�=�~����%�ƿ ؿ[���� �2�u�V� 9�zό�oϰ��ϥ��� ��
�ߟ�=��d�� 9�Ϭ߾�������� ���<�N�1�r��g� ��+ߑ�O���s߅ߗ� ��J���n���c����� ����������4�� ���|���#�5�� ��0B%f I����Ug //�;/�b/t/W/ �/{/�/�/�/�/?�/ (??L?^?��f?�? )/?M/�? OC?$OO 5OZO=O~O�OsO�O�O �O�Om?_�?2_�?_ �?z_�_�O�_�_�_�_ �_
oo�_@oRo5ovo �O___�oA_S_e_�o [o<N1r�g ��������o �oJ�\��o}���� ��ڏ������4�� E�j�M�����#�5�֟ �k�����0�B���f� I��������ү���� ٯ�,���M��t��� I����ο���� (��L�^�Aςϔ�w� ��;���_� ߃����� �Zߝ�~ߐ�sߴߗ� ������� ��D��� )��`�V�������������8�7�I�^�=�H���2k�  �����{����������`����FXj g��C(  @@  �A�Ӈ@�{�A   ?��?р� � g�@��f�fC�!�	 B�p� �  F?1����@�l#��   B� B_�  C��� �`!�H�f�� �A 5�L���� ������ � �A� ��� �$D�CSS_CNST�CY 2P���  md����//4/B/ T/f/|/�/�/�/�/�/��/�/??,?>?�D�EVICE 2QB�#�5"�&�T? _��?�?�?�?�?OO (OUOLO^O�O�O�O�O �O�O�O	__-_�F��HNDGD R��$�Cz��LS 2S��_�_ �_�_�_�_oo:_��PARAM T��bT��Q�2��RBT 2V�� 8 
 < �?} � ���� �E��R�8�l�a�Ĺ0�W  �eB�\�o�f���Cpĉ%.w#��o�f>P�K0�����q$��n� ��f����|�b�u���Fc Rj� ��]�4�F�e�j��|����IC��D�jPC�$Z��@����A,��4��u@�X@���^@w���J��B�%���C4�C3:^oC4��A�����8�-B�{B��A�����&�l��C��C3�JC4�jC3��d� �+�3 Dff 2�A PЩ��K@�d�����ן� ����l�C�U���y� ��������ӯ ���	� V�-�?�Q�c�u���Կ ����
�ϗ�4�F�1� j�Uώ�yϲϝ����� ğ��ڿ��g� >�Pߝ�t߆ߘߪ߼� ������Q�(�:�L� ^�p��������� �� �M���q�\����� ������������� .�#�DV�z� ������
W .@�dv��� �/��A//*/I/ �/�/�/�/�/�/�/ �/+??O?*X/j/�? R/�?�?�?�?�?O�? �?KO"O4OFOXOjO|O �O�O�O�O�O�O�O_ _0_}_T_f_�_�_@? �_�_o�_1ooUo@o Ro�of?�_�_�o�o�o 	�o�o(:� ^p������ �;��$�q�H�Z�l� ~������jo��%�� I�4�m�X���|���ǟ �oЏ�����E�� .�M�R�d�v�ï���� ��Я����*�w� N�`�����������̿ ޿+Ϧ�O�:�_υ�p� �ϔ��ϸ���̟ޟ� ����"�4߁�X�j߷� �ߠ߲�������5�� �k�B�T�f�x��� �����������g� �ϋ�v������������	��-:	�$DC�SS_SLAVE W���[��D
_4�D  [pAR�_MENU X[ "����6��@R@�SHOW 2Y[ � /?� ������/"/(F/X/j/ ��/� �/�/�/�/�/?4/1? C?U?|/v?�/�?�?�? �?�?�??O-O?Of? `O�?�O�O�O�O�O�O O__)_POJ_tOq_ �_�_�_�_�_�O�_o o:_4o^_[omoo�o �o�o�_�o�o�o$o HoEWi{���o @��,2/�A� S�e�w��������я ����+�=�O�a� s������������ ���'�9�K�]�o��� ������ޟد���� #�5�G�Y���}����� ȯ¿������1� C�j�g�yϋϲ���ֿ ������	��-�T�Q� c�uߜϖ��Ͻ����� ����>�;�M�_�� ��ߧ��������� (��7�I�p�j���� �������������!�3eCFG Z�{������FRA:\s�L}%04d.C�SV@	 }@ m�A �CH� �zd��[�����h�.@R>��JP�n2  AS�RC_OUT -[^h���_C_FSI ?��  �&////X/S/e/ w/�/�/�/�/�/�/�/ ?0?+?=?O?x?s?�? �?�?�?�?�?OOO 'OPOKO]OoO�O�O�O �O�O�O�O�O(_#_5_ G_p_k_}_�_�_�_�_ �_ o�_ooHoCoUo go�o�o�o�o�o�o�o �o -?hcu �������� �@�;�M�_������� ��Џˏݏ���%� 7�`�[�m�������� ǟ�����8�3�E� W���{�����ȯïկ ����/�X�S�e� w������������� �0�+�=�O�x�sυ� ���ϻ�������� '�P�K�]�oߘߓߥ� ����������(�#�5� G�p�k�}������ �� �����H�C�U� g��������������� �� -?hcu ������� @;M_��� �����//%/ 7/`/[/m//�/�/�/ �/�/�/�/?8?3?E? W?�?{?�?�?�?�?�? �?OOO/OXOSOeO wO�O�O�O�O�O�O�O _0_+_=_O_x_s_�_ �_�_�_�_�_ooo 'oPoKo]ooo�o�o�o �o�o�o�o�o(#5 Gpk}���� � ����H�C�U� g���������؏ӏ� �� ��-�?�h�c�u� ��������ϟ���� �@�;�M�_������� ��Я˯ݯ���%��7�`�[�m��$DC�S_C_FSO �?������ P  s�m���߿ڿ���'� "�4�F�o�j�|ώϷ� ������������G� B�T�fߏߊߜ߮��� ��������,�>�g� b�t��������� ����?�:�L�^��� �������������� $6_Zl~� ������7 2DVz��� ���/
//./W/ R/d/v/�/�/�/�/�/��/�/�C_RPI����
?S?|?w?"?���F?�?�?�?�?��SL4?@�?OQOzOuO �O�O�O�O�O�O
__ _)_R_M___q_�_�_ �_�_�_�_�_o*o%o 7oIoromoo�o�o�o �o�o�o!JE Wi������ ��"��/�A�j�e� w���������я���� ��B�=�O�a����� ����ҟ͟ߟ���  O�?DO&�o������� ���ۯ���(�#�5� G�p�k�}�������ſ ׿ �����H�C�U� gϐϋϝϯ������� �� ��-�?�h�c�u� �߽߰߫�������� �@�;�M�_���� ������������%� 7�`�[�m�������� ��������83�<�NOCODE }\�5��;�PRE_CHK �^�;J A J �< �O �5���5 	 < �W��=O) s�_q���� /�'/9//%/o/�/ [/�/�/�/�/�/��/ #?5?�/Y?k?E?w?�? {?�?�?�?�?OO�? +OUO/OAO�O�OwO�O �O�O�O	_�/??_Q_ �O]_�_a_s_�_�_�_ �_o�_o;oo'oqo �o]o�o�o�o�o�o�o �o%7[m'_U �������!� ��W�i�C�����y� ÏՏ��������A� S�-�w���q���џ k������=��)� s���_�������ǯ� ˯ݯ'�9��]�o�I� {�������ۿ���� #����Y�k�EϏϡ� {ϭ��ϱ������� C�U�/�aߋ�e�w��� �߭���	�ÿ��?�Q� +�u��a����� �����)�;��_�q� K�]������������� %�[m� �}����! �EW1c�gy ����/�/A/ 7Iw/�/#/�/�/�/ �/�/?�/+?=??I? s?M?_?�?�?�?�?�? �?�?'OOO]OoOIO �O�O_/�O�O�O�O_ #_�OG_Y_3_E_�_�_ {_�_�_�_�_o�_�_ CoUo/oyo�oeo�o�o �O�o�o	�o-? KuOa���� ���)���_�q� K���������ݏ�o�o �%���1�[�5�G��� ��}�ǟٟ����� ��E�W�1�{���g��� ï��������/�A� ��)�w���c������� ���Ͽ�+�=��a� s�Mϗϩσϕ����� ���'��K�]�S�E� �ߥ�?����ߵ���� ����G�Y�3�}��i� �����������1� C��O�y�o߁߯��� [���������-? cuO����� ��)5_9 K�������� /%/�I/[/5//�/ k/}/�/�/�/�/?�/ 3?E??1?{?�?g?�? �?�?�?�?��?/OAO �?eOwOQO�O�O�O�O �O�O�O_+__7_a_ ;_M_�_�_�_�_�_�_ �_oOOKo]o�_io �omoo�o�o�o�o �oG!3}�i �������1� C��g�y�3oa����� �����я�-��� c�u�O�������ϟ� ��͟�)��M�_�9� ������}�˯ݯw�� ���I�#�5���� k���ǿ��ӿ��׿� 3�E��i�{�Uχϱ� �������ϓ��/�	� �e�w�Qߛ߭߇߹� �߽����+��O�a� ;�m��q������� ������K�]�7��� ��m����������� ��5G!k}Wi ������1 '�gy��� ����/-//Q/ c/=/o/�/s/�/�/�/ �/??�/#?M?CU �?�?/?�?�?�?�?O O�?7OIO#OUOOYO kO�O�O�O�O�O�O	_�3___i_{_����$DCS_SGN� _k5��%)��1�8-JUL-24 12:10 ]S�05-MAR>�Q00:41�P�P��R Xza�E�RehXe�U�Q�R�Y�P�Q�R�B,�Þ����E��_�Po�����5��X���K�_U�THO�W `k5� �Q�UVE�RSION ��V�`�V4.�5.8�Y�PEFLOGIC 1aui?�  	\Pf�p0�ip0�n�bPRO�G_ENB  ��T�c�P	sULSOE  �e!u�b_ACCLIM4v��#sdHsW?RSTJNT4w�a;��TEMO|�Q�%q�b�pINIT �b�jg:�`�tOPT_SL ?	k6��r
 	R5�75�S�p74�y6Z�x7�w50�1��2�t�hG��g�tTO�  �}#o���fV.�pDEX4wd�b�P���PATH �A�jA\ 80�72024\ U�ME INFORMAT�`\����c�HCP_CLNT�ID ?�f�c ��h�UR��bIA�G_GRP 2gvk5a��R	 @�  ��ff?aG���<�Z��B�  ȟ�\�ő�ΐ�ߞ@c����!�7@�z��@^�@
��!�Ymp3m�29 8901234567E��ws0w� ����Rd�`h�}��Va��QB4�����X �U�xͣ a�_�k6���>�k6 Ѡc>������-�ǿ8Q�c�u��\�Կ Ϩ���T�޿�Ϝ� ��8϶���nπϒ�,� >���b�t���l�xߺ� Dߪ�������8�J� (�Z��
��f����� �������4�q2c�d�x!� Ѹ�?��x��@`������5!=���4V������A�P��@����Z��?����������8��F�=q�=b���=�E1>�J��>�n�>���H��<�o D
�SsT�\N���Q�Cp  <(�U.�R 4������-��YA@�R?�� �@���i8� F�V|^��D��>J���bN<�����G�����@���$"��?��0!@f�f�!6 M!33ܳX"(�ø�C��� t"I�CH��)C.dB؃���΢�/�!�,' 6p�/��͐�%B�P�%Xd.[ 1B���7�/=?O?B XT�G�����ҟ?��]���?\��?�����J>��~�.I�d���CD23D4�3�P(��� Q?�?�?�?�(�?B�R9�9Ca~�������;;���?UO@OyOdO�O��O�O�OR39����;�ܺ����<���;D�=�U:�oUn��CT_CONFI/G h���s�T�eg�ez�STBF_TTS4w�
!yhS�`4s�Q{V�h`MAUop�bM_SW_CF<Pi���  �lOCVI�EW�Pj�]Ñ��g�!o3oEoWoio{o MRo�o�o�o�o�o�o �o"4FXj| �������� 0�B�T�f�x������ ��ҏ������,�>� P�b�t�����'���Ο �������:�L�^��p�����$\PM�R�k�]RSͧШ
 �έ����SCH� 2r�[
|�Schedul'e 18k oRQ`
R4��`��*3ϥ���]�R;��MQ>L�ͯ���ܿ����˿ $����l�7�I�[� ��ϑϣ��������� D��!�3ߌ�W�i�{�8�ߟ߱�	 l����`��PST�`	�� R9Dz.����#�5�G� Y�k�}�������� ������1�C�U�g� y��������������� 	-?Qcu� ������P);M�NR5=�� ������//)/;/M/_/q*	���/�/ �/��I VB�T�?x� ��K?�߸�:?�?^?p? �?�?�?�?�?#O�? O OkO6OHOZO�O~O�O �O�O�O�O�OC__ _ 2_�_V_ �r��� �`�_�_�_�_
oo .o@oRodovo�o�o�o �o�o�o�o*< N`r����� ����&�8�J�\� n���������ȏڏ� ���~/|/����ԟ ���
���/L�^�p��/�"%�21��/?� )?{_��_i_�`�+� =�O���s�����𿻿 Ϳ߿8���'π�K� ]�o��ϓϥϷ���� ����X�#߱_#�5�G� Y�k���ߡ߳����� ������1�C�U�g� y������������ 	��-�?�Q�c�u��� ������������ );M_q��� ��}�/�Yk}� ����1�C�/+/ =/���/˯�/�A��/ e�/߱/
?�/�/�/R? ?/?A?�?e?w?�?�? �?�?�?*O�?OOrO =OOOaO�O�O�O�O_ �Ow���1�_ 9_K_]_o_�_�_�_�_ �_�_�_joo#o5oGo Yo�o}o�o�o�o�oB �o�o1�Ug y������� 	���-�?�Q�c�u�� U��'�9�K�]�o� ����	/ß՟�Q/����3��o/�/^��/�O ��_�O��ܯ����˯ $����l�7�I�[� ���������ǿٿ� D��!�3ό�W�i�{� �ϟ�-_����ÏՏ� ����/�A�S�e�w� �ߛ߭߿�������� �+�=�O�a�s��� �����������'� 9�K�]�o��������� ��������#5G �������/ AS�������� i/G�/k���>/�ϫ� -/�/Q/c/u/�/�/�/ �/?�/�/?^?)?;? M?�?q?�?�?�?�?�? �?6OOO%O~OIO�� ew���_�O�O �O�O�Oz_!_3_E_W_ i_�_�_�_�_�_�_Ro �_oo/oAo�oeowo �o�o�o*�o�o�o �=Oas�� �����n��o ������Ǐُ������?�Q�c���%�4 )���ڟ!/sO��O aO��X�#�5�G���k� }���诳�ůׯ0��� ��x�C�U�g����� �����ӿ���P�� �O�-�?�Q�c�	��� �ϫϽ��������� )�;�M�_�q߃ߕߧ� ����������%�7� I�[�m������� �������!�3�E�W� i�{���������u�'� Qcu����� )�;�#5���ß ��9Ϻ]�'ϩ/ ���J//'/9/�/ ]/o/�/�/�/�/�/"? �/�/?j?5?G?Y?�? }?�?�?�?�?o����� )�O1OCOUOgO yO�O�O�O�O�O�Ob_ 	__-_?_Q_�_u_�_ �_�_�_:o�_�_oo )o�oMo_oqo�o�o �o�o�o�o~%7 I[m�M��� 1�C�U�g�y����� ͏ߏI����5��g yV���?��O�?{� ԟ����ß����� d�/�A�S���w����� ����ѯ�<���+� ��O�a�s�̿��%O� �������'� 9�K�]�oρϓϥϷ� ���������#�5�G� Y�k�}ߏߡ߳����� ������1�C�U�g� y������������ 	��-�?�������� ��'9K���� �����a?� c� ��6ٿ��%~I[ m����/�� �V/!/3/E/�/i/{/ �/�/�/�/�/.?�/? ?v?A?�]�o����� ��O�?�?�?�?�?rO O+O=OOOaO�O�O�O �O�O�OJ_�O__'_ 9_�_]_o_�_�_�_"o �_�_�_�_o�o5oGo Yoko}o�o�o�o�o�o �of��g���� ����}7�I�[����6!���ҏ k?��?Y?��P�� -�?���c�u������� ��ϟ(����p�;� M�_��������� �˯ ݯ�H���?%7 I[�������ǿ ٿ����!�3�E�W� i�{ύϟϱ������� ����/�A�S�e�w� �ߛ߭߿�������� �+�=�O�a�s��� ���m�I�[�m�� ��������!�3�	 -{����|ߏ1�� U�������B 1�Ugy� ���/��	/b/ -/?/Q/�/u/�/�/�/ �/g��������!��? )?;?M?_?q?�?�?�? �?�?�?ZOOO%O7O IO�OmOO�O�O�O2_ �O�O�O_!_�_E_W_ i_{_�_
o�_�_�_�_ �_voo/oAoSoeo�o E���);M_ q������A����7��_qN���/ ��?�/s�̏������ �ߏ��\�'�9�K� ��o�����쟷�ɟ۟ 4����#�|�G�Y�k� į��?�o�o�o�o�o }o����1�C�U�g� y���������ӿ��� 	��-�?�Q�c�uχ� �ϫϽ��������� )�;�M�_�q߃ߕߧ� ����������%�7� �o����������� 1�C���������� Y7���[���.ѯ�� vASe��� ����N+ =�as���� �&/�//n/9/� U�g�y����/�/�/ �/�/�/j??#?5?G? Y?�?}?�?�?�?�?BO �?�?OO1O�OUOgO yO�O�O_�O�O�O�O 	_�_-_?_Q_c_u_�_ �_�_�_�_�_^o��_� �o�o�o�o�o�o�o�o�u�/AS����8 ������c/ ��/ Q/�H��%�7���[� m��؏����Ǐ �� ���h�3�E�W���{� ������ß՟�@�� �/oo/oAoSo�_w� ��������ѯ���� �+�=�O�a�s����� ����Ϳ߿���'� 9�K�]�oρϓϥϷ� ���������#�5�G� Y�k�}ߏߡ߳�eo A�S�e�w����� +��%�s��� t��)���M������ ������:)� M_q���� ��Z%7I� m���_����� ����z/!/3/E/W/ i/�/�/�/�/�/�/R? �/??/?A?�?e?w? �?�?�?*O�?�?�?O O�O=OOOaOsO�O_ �O�O�O�O�On__'_ 9_K_]_�_=����_o !o3oEoWoio{o��o �o�o9��p9�W� i�F���|/�k �������� T��1�C���g�y��� 䏯���ӏ,���	�� t�?�Q�c�����/�_ �_�_�_�_u_��� )�;�M�_�q������� ��˯ݯ���%�7� I�[�m��������ǿ ٿ����!�3�E�W� i�{ύϟϱ������� ����/��_�o���� ������)�;�o�o }����oQ�/��S ��&�ɟ���n�9�K� ]��������������� ��F#5�Yk }������ f1۟M�_�q߃� ��������b/ 	//-/?/Q/�/u/�/ �/�/�/:?�/�/?? )?�?M?_?q?�?�?O �?�?�?�?O~O%O7O IO[OmO�O�O�O�O�O �OV_��W�y_�_�_�_ �_�_�_�_m�'o9oKo4���hv10w ��o�T�oxB�o 9(�L^p ������� � Y�$�6�H���l�~��� 鏴�Ə؏1����� _ _.�D_���Oz��� ����-�ԟ���
�� ��@�R�d�v������ ��Я���q��*�<� N�`�ݿ��������̿ I����&�8ϵ�\� nπϒϤ�!�h_oD� V�h�zߌߞ߰���o ����do��o�ow� �oh��P������� ��������,�>�P� b�t������������� ��(:L^p ����b������� 
����$6HZl ~������� / /2/D/V/h/z/�/ �/�/�/�/�/�/
?? .?@?R?d?v?�?�?�? �?�?�?�?OO*O<O NO`O.����O __$_ 6_H_Z_l_��$�_�_�*�<��$DRC_�CFG sE��!L�o�J oKo:ooo^o�o�o�o���PSBL_FA?ULT t	j�e��dGPMSK  ��d�g�PTDIA�G uE��Q�P����UD1: 67�89012345�Ar�5q\��P  �o������ ��!�3�E�W�i�{� ���oY�4s��@�Cm|��eTRECP,z
:t,�Sw/�kh� z�������ԟ��� 
��.�@�R�d�v���௏��ӏЯ�gUMP_OPTION�`��n�TRb�c�i��PMES�	�Y�_TEMP  ?È�3B�� _���A\�I�UNIT��g_�vYN_BR/K v	�(r��?EDITOR����8���_�ENT �1w	i�@,&�ROS2  OR�r����J&PRO�VA��2�&	T�RANSP"�4�&DE�c{�
Χo�������������� �5��Y�@�}ߏ�v� �ߚ����������1� �*�g�N��r���� ������	���?�&����MGDI_ST�Ar��_�� ��N�C_INFO 1�x��������`3����~�f�1y�� ������� �E d��M_q�� �����% 7I[m��� ����//"): "/H/Z/l/~/�/�/�/ �/�/�/�/? ?2?D? V?h?z?�?�?�?**� �?�?OO1/;OMO_O qO�O�O�O�O�O�O�O __%_7_I_[_m__ �_�_�_�?�_�_�_o )O3oEoWoio{o�o�o �o�o�o�o�o/ ASew����_ ����!o�=�O� a�s���������͏ߏ ���'�9�K�]�o� ��������۟��� ��+�5�G�Y�k�}��� ����ůׯ����� 1�C�U�g�y������� ɟӿ���	�#�-�?� Q�c�uχϙϫϽ��� ������)�;�M�_� q߃ߕߧ��������� ��%�7�I�[�m�� ������������� !�3�E�W�i�{����� �����������/ ASew���� ���+=O as������� �'/9/K/]/o/ �/�/�/�/�/�/�/�/ ?#?5?G?Y?k?}?�? ���?�?�?�?/O 1OCOUOgOyO�O�O�O �O�O�O�O	__-_?_ Q_c_u_�_O�?�_�_ �_�_Oo)o;oMo_o qo�o�o�o�o�o�o�o %7I[m ��_����o� !�3�E�W�i�{����� ��ÏՏ�����/� A�S�e�w�������� џ����+�=�O� a�s���������ͯ߯ ���'�9�K�]�o� ��������ɿۿ��� �#�5�G�Y�k�}Ϗ� �ϳ����������� 1�C�U�g�yߓ����� ��������	��-�?� Q�c�u������� ������)�;�M�_� q����ߧ��������� %7I[m ������� !3EWi{��� ������//// A/S/e/w/�/�/�/�/ �/�/�/??+?=?O? a?s?�?�?�?�?� �OO'O9OKO]OoO �O�O�O�O�O�O�O�O _#_5_G_Y_k_�?�? �_�_�_�_�?�_oo 1oCoUogoyo�o�o�o �o�o�o�o	-? Qc�_�_���� �_���)�;�M�_� q���������ˏݏ� ��%�7�I�[�m�� ������ǟ����� !�3�E�W�i�{����� ��ïկ�����/� A�S�e��m������� ٟϿ����+�=�O� a�sυϗϩϻ����� ����'�9�K�]�w� ���ߥ߷�m������ �#�5�G�Y�k�}�� ������������� 1�C�U�o߁ߋ����� ��������	-? Qcu����� ��);M_ y��������� //%/7/I/[/m// �/�/�/�/�/�/�/? !?3?E?W?q{?�?�? �?��?�?�?OO/O AOSOeOwO�O�O�O�O �O�O�O__+_=_O_ i?[_�_�_�_�?�?�_ �_oo'o9oKo]ooo �o�o�o�o�o�o�o�o #5Ga_s_}� ���_����� 1�C�U�g�y������� ��ӏ���	��-�?� �ku��������ϟ ����)�;�M�_� q���������˯ݯ� ��%�7�I�c�m�� ������ǿٿ���� !�3�E�W�i�{ύϟ� ������������/� A�[�I�w߉ߛߵ��� ��������+�=�O� a�s��������������'�9�S� ��$ENETMOD�E 1z����  c��c�^Հ���b�OATCFG {��/������C���DATA �1|o����**��1C$Uddd��������k�� ��Zl~����7I�//,/�P/�����/�/ �/�/?/�/��o/�/�.?@?R?d?�/�?�� ??�?�?�? Ow?$O���?�?fOxO�O�O�O�OZ�RPOST�_LO��~��^�
���	__-_?_�BROoR_PR�@%o��%]�x_G_R_TA�BLE  o�����_�_�_�WSRSE�V_NUM ~��4�y�`�A_�AUTO_ENB�  ��w��D_N�O-a o����b  *�p`�Jp`�p`�p`#`+o`��o�o�oIdFLTR5oGfHISc2@m_ALM 1�o�� �g%pl]�+ �oI[m���o�_bO`  o��na���zb�TCP_�VER !o�!�p_�$EXT�@_7REQ�f�@i:��SIZC�5�STK�`�^e�7�TOoL  `�Dz�b��A 5�_BW�D�p���fɁ��DI�� ����G��<�ϊSTEPߏ�|b��OP_DO���`�FDR_GRP� 1�o��ad 	������q�s�V���'�N"����l��T� �����q�Ɵ ם������	�B�-�� ? �����̾2�\=�ʾ�z?T���P����ï^��Β@A�Z}@1�>ҿ�Z=(��Ǫ
? ML�`��l�ǯv��ȯ��W�xB�{�f�A@  ��O@S33��`�@�����_����q�F@� �ռq�G�  �8�Fg�fC�8RD�ؽ?�f�a�׾�6�X����87�5t��5����5`+�ؽ���\���JY���Ǔ���7�p�m�KFE�ATURE ����ɀ��L�R HandlingTool ��`�Engli�sh Dicti�onary�4Dw St��ard���Analog �I/O6�?�gle� ShiftR�u�to Softw�are Upda�tew�matic Backup����ground �Edit���Ca�meraM�FQ�C�ommon ca?lib UI�����n����Monit�or �tr �Re�liabf��DH�CP���Data Acquis�~8�iagnos���J�R�isplay~��Licens6��<�ocument? Viewe�:��ual Chec�k Safety����hancedh�����s��Fr����xt. DIO� �fi���en]d��Err�L��8��s7�rH�'� ����FCTN M�enu��v6��T�P Iny�fac<���GigE�������p Mask �Exc��g�HT���Proxy S�v����igh-S;pe��Ski�������+�mmunicn��ons2ur���y�M�Nѳ�conn�ect 2inc=r��stru�g
�� e����J���K�AREL Cmd7. L��ua����Run-Ti�E�nv�z�el +:��s��S/Wע������N�Book(System)�MACROs,)?/Offsem�LaH+���K�QMR�D��M��| *�l���MechStop"t� l�LiI�i���x��JТ�{od>g�witch/��{�.q,+Optm�>/� fi��g�_Lulti-T������PCM f�un��)a�ti�z�(�'oi�RegeiArM �&ri���F�+6K�Num �Sel�'9� Adju= ">O1i�`=tatu1x?����RDM Robo}t�scove��5ea� �Fre�q AnlyMRem�+�n-״5�2Servo+� �?SNPX b	n�;SN��Cli��7Nj�Libr�WO��Q �i@#Fo&t���ssag�%�D�p 0�d9��p/I���E�MILIB�O�BP� Firm���NPΗ�Acc����TPsTXG�Delnd��O�A��`�Morq}ug�imula�4��tVu  Pa�N��4�:#& ev.̰E��ri��L_USR EVNT�_�`nexcept����0n�� e�S�VEC��rH?�Vh�eb_veiKpkSJ@S9CFU�oSGE�o�e�UI9�Web Pl�6�nA_t �����n�ZDT Ap�plF�WqEOA�T�A���iPB�a|PI� Grid�1���}|iR\b.�-��v{�}o��RX-�10iA/L�A�ll Smoot�h-��s�S���Pr�ityAvoidM�s/�t�P?���bV0o���!��ycf�`�0�P��;�CS�� . c�⼈Jo 1� ф׏$҂�����M�|��c�abo��4��main N�A.8�yp y� �ifi����PMC����RL�P�
y&��av����p��bc~��MI Dev�� (+AE�y�d�1/��ַS��"��1�0iC�rt(�e1n��4��ni+�x�!���'sswo4���ROS Eth��P��eMw�4��9LX� b���E<�UapN0A�E3�t �����Wr0 dow�n-al�Puero DN��V ��z�
v��vK4��8�64MB� DRAM4���F�RO��}�X�� F!l  �0`�� r�2�os�n�Ce8�N���#shD�P�b�c]+_Ų��p�Vt�tyf�s 92����ᯧ��2V _���́/s���d���0k�O�� 2��a�|�por*�EMAILB{~�Q���MK���0B.�q��T1��FChe��Fs��Hel�u�޿3�Typ��FC h��*`SLFor0��(�r�lu �4<2�LCMGRH_NOPG j�}R�z�z/�1reP0)�Ne�tFr)г���o �m�0�0c���tOPOC-UA��3�T1�Ȕ A���S�p��cr�ꀲ+lu�@ AP �e����!(7( �3�t�:�Qp�PSyn�.(RSS)�6q?uires �@'���3iE�tN���es�t�EIMPLE @��f"G��LM#FS��e�Btex�T���!HplQ3b�_CPP ExO�?+��`x�Tea  tY���VɠF��ru�&(�!S���QСxۑ��@�fUI�Fƒoni��ust'dpn�[�t��r� �����+/"/4/ F/X/�/|/�/�/�/�/ �/�/�/'??0?B?T? �?x?�?�?�?�?�?�? �?#OO,O>OPO}OtO �O�O�O�O�O�O�O_ _(_:_L_y_p_�_�_ �_�_�_�_�_oo$o 6oHouolo~o�o�o�o �o�o�o 2D qhz����� ��
��.�@�m�d� v�������ُЏ�� ��*�<�i�`�r��� ����՟̟ޟ��� &�8�e�\�n������� ѯȯگ����"�4� a�X�j�������ͿĿ ֿ�����0�]�T� fϓϊϜ��������� ����,�Y�P�bߏ� �ߘ��߼�������� �(�U�L�^���� ��������� ��$� Q�H�Z���~������� �������� MD V�z����� ��
I@R v������� //E/</N/{/r/�/ �/�/�/�/�/�/?? A?8?J?w?n?�?�?�? �?�?�?�?�?O=O4O FOsOjO|O�O�O�O�O �O�O�O_9_0_B_o_ f_x_�_�_�_�_�_�_ �_o5o,o>okoboto �o�o�o�o�o�o�o 1(:g^p�� ����� �-�$� 6�c�Z�l�������Ϗ Ə؏���)� �2�_� V�h�������˟ԟ ���%��.�[�R�d� ������ǯ��Я��� !��*�W�N�`����� ��ÿ��̿޿��� &�S�J�\ωπϒϿ� ����������"�O� F�X߅�|ߎ߻߲��� �������K�B�T� ��x���������� ���G�>�P�}�t� ������������ C:Lyp�� ����	 ? 6Hul~��� ��/�/;/2/D/ q/h/z/�/�/�/�/�/ ?�/
?7?.?@?m?d? v?�?�?�?�?�?�?�? O3O*O<OiO`OrO�O�O�O�O�F  ?H551�C�A�2�FR782�G5�0�EJ614�EAwTUPV545X�6�EVCAM�EC�UIFW28[VN�REV52NVR6�3WSCH�ELI�C~VDOCV�VC�SUV869W0^*VEIOCW4V�R69NVESET�7WMWJ7MWR68��FMASK�EPR�XYgX7�FOCOBh37XV`X3Vf[J6X53�VH�h�LCH>fOPLGz7W0nfMHCR?f�S�gMAT~VMC�S6X0g55*VMgDSW#wagOPagGMPRbf�P�h0VPCMfW5iw`*Vl�`�g51BW51�x�0BVPRSg69�VfFRDZVFRE�QVMCN�F93�VSNBA�W�gSHLB�M)��Px�2VHTC6VTMsILX�VTPA�VoTPTX[�EL�v��`�W8WP�FJ9�5rVTUTbfUE�VfUEC>fUF]RZVVCC��O�fwVIPf�CSC���CSG~V�PI�EW�EB6VHTT6VRa6�X��3P>�CGU�{IG=�IPGS���RCf�DGagH7X�w�`W51�X6nh�0rVK�nh5NV�PJ�x�x6rWL)�J7v!�R7�gS50W�̘J64�VR55`nf�rV�P�w76hU7�FS�Z4��5ɧ�R6�gR9٘79bzh4rV��VfWN	w�R8!wR76BW7]6VfD06*VFL�wRTS�CRDfwCRXbfCLIRx�AWCMS�V��6VS�TYf�6!wCTO�6V�P�W7�W�P�N9N��VfORS�f/`�VFCB�VFCFv�wCH6VFCRf�FCI��FC�gJ����gM�gPG�M��xR58*VNET�fVNOM�VCp�VO�Pa�SEND?fAP>�PLU�f�P��]7�VCPR�wL��S�C�Y67VfE�TS�Ǡ��Pr�CP�~VTEq�S6]�T�OA.vTRA>fI�N�wIHY�IPN f��H������%�7� I�[�m������� �������!�3�E�W� i�{������������� ��/ASew ������� +=Oas�� �����//'/ 9/K/]/o/�/�/�/�/ �/�/�/�/?#?5?G? Y?k?}?�?�?�?�?�? �?�?OO1OCOUOgO yO�O�O�O�O�O�O�O 	__-_?_Q_c_u_�_ �_�_�_�_�_�_oo )o;oMo_oqo�o�o�o �o�o�o�o%7 I[m���� ����!�3�E�W� i�{�������ÏՏ� ����/�A�S�e�w� ��������џ���� �+�=�O�a�s����� ����ͯ߯���'� 9�K�]�o��������� ɿۿ����#�5�G� Y�k�}Ϗϡϳ������  H5�5������2��R7�82��50��J6;14��ATU��5��545/�6��VC{AM��CUIF/ۻ28�NRE�5�2n�R63�SC�H��LIC��DO�CV��CSU�8�69/�0>�EIOuC��4�R69n��ESETO�m�J7�m�R68�MAS�K��PRXY��7.��OCOo�3O�ڴ{�.�3��J6-�5u3�H�LCH��OPLGO�0��M�HCR��Sm�MA]T��MCSN�0~�{55>�MDSW��v��OP��MPR��t���0.�PCM���5={�>�{��51�^�51~0^�PR�Sn�69��FRD�~�FREQ�MC�N��93.�SNByA���SHLB�M=����2.�HT=CN�TMIL���TPA>�TPTXFEL�
{��8����J95��TU�T��UEVn�UE�C��UFR~�VCuCN,O��VIP�wCSC�CSG�ں�I��WEBN�HTTN�R6���Kж�*CG�+IG�+I�PGS:RC�D�G��H7�+��51N�6��0��k��I5n��J���6��mL=J7�;R7=��S50�l<J64�R55��[@��[�Vn76~�7�S�޵4�5�KR6}�R-9}<79��4�ګ@���WN��R8��R�76^�76��D0u6>�Fl\RTSwCRDn�CRX���CLI]�CMS�>��PN�STY�6���CTON��>�7��О;NNNm��O�RS����.�FCBn>�FCF�CHN�wFCRn�FCI.:KFC��J0��M���PG�:M�R58�>�NET��NOM�>� �OP�kSE�ND��AP�*PL�Un��nL7�CPUR�L]+S|lC�;67��ETS~{�\l+��CP��TE�[�S6-KTOA��T�RA��IN�IH}IPN���Տ� ����/�A�S�e�w� ��������џ���� �+�=�O�a�s����� ����ͯ߯���'� 9�K�]�o��������� ɿۿ����#�5�G� Y�k�}Ϗϡϳ����� ������1�C�U�g� yߋߝ߯��������� 	��-�?�Q�c�u�� ������������ )�;�M�_�q������� ��������%7 I[m���� ���!3EW i{������ �////A/S/e/w/ �/�/�/�/�/�/�/? ?+?=?O?a?s?�?�? �?�?�?�?�?OO'O 9OKO]OoO�O�O�O�O �O�O�O�O_#_5_G_ Y_k_}_�_�_�_�_�_ �_�_oo1oCoUogo yo�o�o�o�o�o�o�o 	-?Qcu� �������� )�;�M�_�q������� ��ˏݏ���%�7� I�[�m��������ǟ ٟ����!�3�E�W� i�{�������ïկ� ����/�A�S�e�w� ��������ѿ���� �+�=�O�a�sυϗ�Щϻ��������STD��LANG����(�:�L� ^�p߂ߔߦ߸����� �� ��$�6�H�Z�l� ~������������ � �2�D�V�h�z��� ������������
 .@Rdv��� ����*<�N`r���R{BT�OPTN� ��//%/7/I/[/ m//�/�/�/�/�/�/��/?!?3?DPN�Q?c?u?�?�?�? �?�?�?�?OO)O;O MO_OqO�O�O�O�O�O �O�O__%_7_I_[_@m__�_�_�_�_�� �_�_	oo-o?oQoco uo�o�o�o�o�o�o�o );M_q� �������� %�7�I�[�m������ ��Ǐُ����!�3� E�W�i�{�������ß ՟�����/�A�S� e�w���������ѯ� ����+�=�O�a�s� ��������Ϳ߿�� �'�9�K�]�oρϓ� �Ϸ����������#� 5�G�Y�k�}ߏߡ߳� ����������1�C� U�g�y�������� ����	��-�?�Q�c� u��������������� );M_q� ������ %7I[m�� �����/!/3/ E/W/i/{/�/�/�/�/ �/�/�/??/?A?S? e?w?�?�?�?�?�?�?��?OO+O=OOOaH��aOO�O�O�O�O�J�99�E�$FEA�T_ADD ?	����
QP  	�H_-_ ?_Q_c_u_�_�_�_�_ �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o �o%7I[m ������� �!�3�E�W�i�{��� ����ÏՏ����� /�A�S�e�w������� ��џ�����+�=� O�a�s���������ͯ ߯���'�9�K�]� o���������ɿۿ� ���#�5�G�Y�k�}� �ϡϳ���������� �1�C�U�g�yߋߝ� ����������	��-� ?�Q�c�u����� ��������)�;�M� _�q������������� ��%7I[m ���������DDEMO �~
Y   �H D:Lyp��� ����//?/6/ H/u/l/~/�/�/�/�/ �/�/??;?2?D?q? h?z?�?�?�?�?�?�?  O
O7O.O@OmOdOvO �O�O�O�O�O�O�O_ 3_*_<_i_`_r_�_�_ �_�_�_�_�_o/o&o 8oeo\ono�o�o�o�o �o�o�o�o+"4a Xj������ ��'��0�]�T�f� ������ɏ��ҏ��� #��,�Y�P�b����� ��ş��Ο���� (�U�L�^��������� ��ʯ����$�Q� H�Z���~�������ƿ ���� �M�D�V� ��zόϹϰ������� �
��I�@�R��v� �ߵ߬߾������� �E�<�N�{�r��� ����������A� 8�J�w�n��������� ������=4F sj|����� �90Bof x������� /5/,/>/k/b/t/�/ �/�/�/�/�/�/?1? (?:?g?^?p?�?�?�? �?�?�?�? O-O$O6O cOZOlO�O�O�O�O�O �O�O�O)_ _2___V_ h_�_�_�_�_�_�_�_ �_%oo.o[oRodo�o �o�o�o�o�o�o�o! *WN`��� �������&� S�J�\����������� �ڏ���"�O�F� X���|�������ߟ֟ ����K�B�T��� x�������ۯү�� ��G�>�P�}�t��� ����׿ο���� C�:�L�y�pςϜϦ� ������	� ��?�6� H�u�l�~ߘߢ����� ������;�2�D�q� h�z���������� ��
�7�.�@�m�d�v� �������������� 3*<i`r�� �����/& 8e\n���� ����+/"/4/a/ X/j/�/�/�/�/�/�/ �/�/'??0?]?T?f? �?�?�?�?�?�?�?�? #OO,OYOPObO|O�O �O�O�O�O�O�O__ (_U_L_^_x_�_�_�_ �_�_�_�_oo$oQo HoZoto~o�o�o�o�o �o�o MDV pz������ �
��I�@�R�l�v� ������ُЏ��� �E�<�N�h�r����� ��՟̟ޟ���A� 8�J�d�n�������ѯ ȯگ����=�4�F� `�j�������ͿĿֿ ����9�0�B�\�f� �ϊϜ����������� �5�,�>�X�bߏ߆� ���߼��������1� (�:�T�^������ �������� �-�$�6� P�Z���~��������� ������) 2LV �z������ �%.HRv �������!/ /*/D/N/{/r/�/�/ �/�/�/�/�/??&? @?J?w?n?�?�?�?�? �?�?�?OO"O<OFO sOjO|O�O�O�O�O�O �O___8_B_o_f_ x_�_�_�_�_�_�_o oo4o>okoboto�o �o�o�o�o�o 0:g^p��� ���	� ��,�6� c�Z�l�������ϏƏ�؏���(�  �>�P�b�t����� ����Ο�����(� :�L�^�p��������� ʯܯ� ��$�6�H� Z�l�~�������ƿؿ ���� �2�D�V�h� zόϞϰ��������� 
��.�@�R�d�v߈� �߬߾��������� *�<�N�`�r���� ����������&�8� J�\�n����������� ������"4FX j|������ �0BTfx �������/ /,/>/P/b/t/�/�/ �/�/�/�/�/??(? :?L?^?p?�?�?�?�? �?�?�? OO$O6OHO ZOlO~O�O�O�O�O�O �O�O_ _2_D_V_h_ z_�_�_�_�_�_�_�_ 
oo.o@oRodovo�o �o�o�o�o�o�o *<N`r��� ������&�8� J�\�n���������ȏ ڏ����"�4�F�X� j�|�������ğ֟� ����0�B�T�f�x� ��������ү���� �,�>�P�b�t����� ����ο����(� :�L�^�pςϔϦϸ� ������ ��$�6�H� Z�l�~ߐߢߴ����� ����� �2�D�V�h� z������������ 
��.�@�R�d�v��� ������������ *<N`r��������&  '!BT fx������ �//,/>/P/b/t/ �/�/�/�/�/�/�/? ?(?:?L?^?p?�?�? �?�?�?�?�? OO$O 6OHOZOlO~O�O�O�O �O�O�O�O_ _2_D_ V_h_z_�_�_�_�_�_ �_�_
oo.o@oRodo vo�o�o�o�o�o�o�o *<N`r� �������� &�8�J�\�n������� ��ȏڏ����"�4� F�X�j�|�������ğ ֟�����0�B�T� f�x���������ү� ����,�>�P�b�t� ��������ο��� �(�:�L�^�pςϔ� �ϸ������� ��$� 6�H�Z�l�~ߐߢߴ� ��������� �2�D� V�h�z�������� ����
��.�@�R�d� v��������������� *<N`r� ������ &8J\n��� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO �O�O�O�O�O�O�O_ _(_:_L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o�o�o�o �o�o�o�o 2D Vhz����� ��
��.�@�R�d� v���������Џ�� ��*�<�N�`�r��� ������̟ޟ��� &�8�J�\�n������� ��ȯگ����"�4� F�X�j�|�������Ŀ ֿ�����0�B�T� f�xϊϜϮ������� ����,�>�P�b�t� �ߘߪ߼�������� �(�:�L�^�p��� ��������� ��$� 6�H�Z�l�~������� �������� 2D Vhz��������
,0 #FXj|��� ����//0/B/ T/f/x/�/�/�/�/�/ �/�/??,?>?P?b? t?�?�?�?�?�?�?�? OO(O:OLO^OpO�O �O�O�O�O�O�O __ $_6_H_Z_l_~_�_�_ �_�_�_�_�_o o2o DoVohozo�o�o�o�o �o�o�o
.@R dv������ ���*�<�N�`�r� ��������̏ޏ��� �&�8�J�\�n����� ����ȟڟ����"� 4�F�X�j�|������� į֯�����0�B� T�f�x���������ҿ �����,�>�P�b� tφϘϪϼ������� ��(�:�L�^�p߂� �ߦ߸������� �� $�6�H�Z�l�~��� ����������� �2� D�V�h�z��������� ������
.@R dv������ �*<N`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o  $6HZl~�� ������ �2� D�V�h�z��������ԏ���
��.��$�FEAT_DEM�OIN  3���^��4�F�INWDEXS�b��F��ILECOMP ��������a�A���SET�UP2 �������  N �ɑ��_AP2BC�K 1��� G �)/����%�0�4����[�1�� �����:����p�� ��)�;�ʯ_���� $���H�ݿ�~�Ϣ� 7�ƿD�m����� ϵ� ��V���z��!߰�E� ��i�{�
ߟ�.���R� ���߈���A�S��� w����<���`��� ���+���O���\��� ���8�����n��� '9��]����" �F�j��5 �Yk���� T�x//�C/� g/�t/�/,/�/P/�/ �/�/?�/??Q?�/u? ?�?�?:?�?^?�?�?� O)O��אP۟ �2�*.SPB�0O{O %FRH�:\PLUGIN	\eO1��0�O�O�5*.VR�O�O�0* �O(_�2-_Q_��HPCY_�_�0FGR6:mR_�Y=_�_�KTr��_o�U�P��_2iU��_Xo�6d@F�O�o�1	�Swa'o�hqEo�oikSTM�o@�R�P�a&o:y�o^ikH�o� wq.p@��nfGIF� �"u���Y�k�nfJPGq���"u��6�0H�ݏ��FJS�����0��S _ˎ
�JavaScri3ptJ�u�CS����!v��>�̍Cas�cading S�tyle She�etsΟ�0
AR�GNAME.DT���<%p\�ȟ҇��R����DI'SP*��>=����M�_���֯��CLLB.ZI󯮯�`K:\�\�oZ�1�CollaboZ���
PANEL1��o��;���T�҇i�Pendant �Panel޿�8	������ɸ(�S�����ϛ�2����Ǹ�� \�nπϒ� �2'�@߀K�.�[���ߘߛ�3 ����Ǹ��d�v߈ߚ� �3/�H�K�6�c����4����Ǹ�� l�~��� �47�P��K�>�k�����)
�TPEINS.X3ML����:\��t����Custom Toolbar�����PASSWORyD?��>FRS˱�CPassw�ord Config��?�Z� O%�I[� ��D�h��� 3/�W/�P/�//�/ @/�/�/v/?�//?A? �/e?�/�??*?�?N? �?r?�?O�?=O�?aO sOO�O&O�O�O\O�O �O_�O�OK_�Oo_�O h_�_4_�_X_�_�_�_ #o�_GoYo�_}oo�o 0oBo�ofo�o�o�o1 �oU�oy��> ��t	��-��� c���������L�� p�����;�ʏ_�q�  ���$���H�Z��~� ����I�؟m����� ��2�ǯV������!� ��E�ԯ�{�
���.� ��տd������/Ͼ� S��wω�ϭ�<��� `�r�ߖ�+ߺ�$�a� �υ�ߩ߻�J���n�������$FIL�E_DGBCK �1�������� < ��)
SUMMA�RY.DG�U�M�D:M����D�iag Summ�ary���CONSLOG��f�x�������� sole� lo���	TPOACCN�l�%T������TP Accountin3����FR6:IP�KDMP.ZIP�����
�����E�xception���y�MEMCH�ECK����|��%�Memory �Data���)���)�RIPE��v��%�� Packets L2����\[�STAT��� %9S�tatus�V	FTP���/��'�mment �TBD*/�w���)ETHERN�Eo/\m/�/��?EthernB)�?figura9��~!DCSVRF/�///?��  v�erify al�l2?��,�%DIFF'???�?3I8diff�?j7\>� CHG01�?�?��?9O��?aO����92/OO(O�O�?^OpO�23�O�O�OA_� �Oh_�FV�TRNDIAG.�LSm__0_�_���Q Ope�#D ~��nostic���	l)VD;EV�RDAT�_�_x�_�_�Vis�Q?Device�_�[IMG�R$o6o�oz2adImagmon�[UP`ESo~�oFRS:\�R}��Updates ListR����`FLEXEVEN�/�o�o����q UIF E�vE!E�{B�)�CRSENSP)K�o����\��/� CR_L�OR_�PEAKZ���PS�RBWLD.CM�����=r��T&�P�S_ROBOWEyLK/�/:GIG��8��\��GigqE�h��S��SM���J�ߟ�~��/EmailcPya����<<)ёHADOW۟��ҟ�g��Shado�w Change���"C�'�RCMERR_�D�V������CFG E/rrorg`t���� ��XcCMSGLIB�ʯܯ`q�t�4��rpic��)��D)]�ZDଟ˿Z�￪ZD成ad���Ό)���T_�_RP��Կ���B�<��$ �Report'��ݤ7�IRDB�EP�ORF�X�j�|�%�iR�gs����{Nt'�NOTI�/�����}߬Not�ific�"��V��) ���<�����p=���,�v�Y� ��}����B���f� ����1���U�g��� �����>�����t�	 ��-?��c��� (�L���� ;�4q �$� �Z�~/��I/ �m///�/2/�/V/ �/�/�/!?�/E?W?�/ {?
?�?.?@?�?d?�? O�?/O�?SO�?LO�O O�O<O�O�OrO_�O +_�O�Oa_�O�_�_&_ �_J_�_n_�_o�_9o �_]ooo�_�o"o�oFo Xo�o|o#�oG�o k�od�0�T� ����C���y� �����>�ӏb����� ��-���Q���u���� ��:�ϟ^�p����)� ;�ʟ_���|��� H�ݯl�����7�Ư [������ ���ǿV� �z�Ϟ��E�Կi� ���ϟ�.���R���v��������$FIL�E_FRSPRT�  �������7�M�DONLY 1��K��� 
 � �ώ��ϲ��Ͽ��߱� ��0�B���f��ߊ� ��+���O������� ��>���K�t����'� ����]�����(�� L��p��5� Y� �$�HZ �~��C�g �/�2/�V/�c/��/5�VISBCK�i�S�x�*.VD��/�/K FR:\�� ION\DAT�A\�/F"K V�ision VD file	?/Q? c?y/�?q/�?:?�?�? p?O�?)O;O�?_O�? �OO$O�OHO�O�O�O _�O7_�OH_m_�O�_  _�_�_V_�_z_o�_ �_Eo�_io{o6o�o.o �oRo�o�o�o�oA S�ow�*<��1�LUI_CON�FIG �K���!�{ $ �sn�{K�3�E�W�i�0{������|x�ŏ ׏�������@�R� d�v��������П� �����*�<�N�`�r� �������̯ޯ�� ��&�8�J�\�n���� ����ȿڿ�����"� 4�F�X�j�|�Ϡϲ� �������ϑ��0�B� T�f�x�ߜ߮����� ��{����,�>�P�b� �߆��������w� ��(�:�L�^���� ����������s�  $6HZ��~�� ���o� 2 DV�z���� �k�
//./@/� Q/v/�/�/�/�/U/�/ �/??*?<?�/`?r? �?�?�?�?Q?�?�?O O&O8O�?\OnO�O�O �O�OMO�O�O�O_"_ 4_�OX_j_|_�_�_�_ I_�_�_�_oo0o�_ Tofoxo�o�o3o�o�o �o�o�o>Pb t��/���� ���:�L�^�p��� ��+���ʏ܏� �� ��6�H�Z�l�~���'����Ɵ؟�������Robot Speed 10%��I�[�m������ � x�����$F�LUI_DATA ����ա���ǤR�ESULT 3��ե�� �T��/wizar�d/guided�/steps/Expert��5�G� Y�k�}�������ſ׿�����Cont�inue wit�h G�ance ��2�D�V�h�zόϞ�`���������� ���-��ե�0� ����A�ա�	�ps�ςߔߦ߸� ������ ��$�6�H� ���o������� �������#�5�G���@ᢟ�G�)ߋ�M�]��cllb�SelectWorkP� ����'9K]�o����Lig�htwe� ��pie���� 1CUgy���� �y����&�]�rip ��To�olNum/NewFram�;/M/ _/q/�/�/�/�/�/�/<�/�0x0�/? -???Q?c?u?�?�?�?p�?�?�?�?  �����3OM�]�!i�meUS/DST �?�O�O�O�O�O�O�O�__+_=_ �Enabl*/q_�_�_�_ �_�_�_�_oo%o7o
Io���!O�o�oWOiF24tO�o�o�o !3EWi{� L_^_������ /�A�S�e�w�����Zo�lo~o��R���ditor��-�?�Q�c� u���������ϟ���� Touch P�anel � (�recommen�)�4�F�X�j�|� ������į֯�ب�����ɏ+�=����accesp߀����� ��ȿڿ����"�4ϾO�Conn�� to Netw�� wωϛϭϿ������� ��+�=߬�_�?��!����!U��In�troductionF��������#� 5�G�Y�k�}����|� �����������*� <�N�`�r��������pOpߒ�����4���cllb�Loa�dSettingNotHW_l�"W���BTfx���������.0 �'9K ]o�������	O������-/���8��!CenterMan��/�/�/ �/�/�/??(?:?� ^?p?�?�?�?�?�?�? �? OO$O6O�//{O�O�5Q/c/u(� 0�O�O_ _2_D_V_�h_z_�_��EOA�T w/o par�O�_�_�_�_oo�0oBoTofoxo�o�� UO���o�o��+�O&��D/DistanceWf�2DVh z������Q? 
��.�@�R�d�v��� ������Џ�MO_OqO�'���&�oz'Offꏄ�������̟ޟ����&�8�S�1 ;�a�s���������ͯ�߯���'�9��
D����oy���%M� _���ֿ�����0�@B�T�f�xϊ�I�2�� �����������!�3߀E�W�i�{ߍ�L���k���?..��/�@S�peedLimit/Max��4� F�X�j�|��������Z	1�p��� 0�B�T�f�x�������`����������Dz��#A,��guid�ed�afety ��u������ �)�[�N` r������� //&/8/g����oW/��/CURegio ſ�/�/�/�/?"?4?�F?X?j?|?�\UTC+01 ~ �23�?�?�?�?�?OO�+O=OOOaOsO�O��
M"}���/i/�O����/	qimezone5�O _2_D_V_ h_z_�_�_�_�_�_���<(�3:00) �Am��rdam, Berlinb�`Rome, Stockhol`?Vienna�_@o Rodovo�o�o�o�o�o�OM!�ѾүO�O#�/�Oe24�oq� �������� %�<I�[�m������ ��Ǐُ����!�3� J/x���#EWv/curren"� ̟ޟ���&�8�J��\�n�����17-�JUL-24 1�P9 ����ί�� ��(�:�L�^�p��������[���Ͽ�� <����Year��� 0�B�T�f�xϊϜϮ�8������20^� �&�8�J�\�n߀ߒ� �߶��������a����#跿!��Month��s�� ������������'���7/�U�g�y� ��������������	0-���� �mr��A𧻓Day2 ����1C0Ugy��1C�� ����//'/9/@K/]/o/�/@R	_p�/ۿ���Hou� ?+?=?O?a?s?�?�?�?�?�?�1�?�?O "O4OFOXOjO|O�O�O �O�O�O�/S�/_�"�/S�inute�Op_�_�_�_�_�_@�_�_ oo$o;�9+o Qocouo�o�o�o�o�o��o�o)�OR		�_i��.=Ucll�b��SetSpe�edLimit/�wVal.��� ��*�<�N�`�r���?250.0��� ����Џ����*� <�N�`�r���A{uCz  _�����rMod^_�&�8� J�\�n���������ȯ���Do not� Use (Re�commen��) ӯ�"�4�F�X�j�|��������Ŀ־ 
8p"8pϟ]�-\})�/Load�p�tingNotHW_lightֿ sυϗϩϻ������� ��ԯZ=�O�a�s� �ߗߩ߻�������� �'�8q걚� �"�t����abSummar���������� �(�:�L�^�p�/ߔ� ���������� $ 6HZl~=�O���5T#��file�2/cyclep/owerKTm� $6HZl~��x���6HOT� �	//-/?/Q/c/u/��/�/�/�/�/�!����?-\9�/ToolP��/d?v? �?�?�?�?�?�?�?O O��<ONO`OrO�O�O �O�O�O�O�O__&_ ��/A_k_�� 5?�{ (_�_�_�_�_oo&o 8oJo\ono-O�o�o�o �o�o�o�o"4F Xj)_;_M_�����_/����%�7� I�[�m��������Ǐ �o����!�3�E�W� i�{�������ß�����(�/Co�nfigurat�ionCompleti�{������� ïկ�����܏A� S�e�w���������ѿ �����ח����?�iχ�XIntroducM�$ϵ��� �������!�3�E�W� i�(��ߟ߱������� ����/�A�S�e�w���Hϒ��.<gui�ded�tNetMethodx��� ,�>�P�b�t�����������Not cE�e����/A Sew����~�  ���y_�s�file/bac�kup�tdevicX�]o���������/|�F�ront Pan�el USB (UD1)/U/g/y/ �/�/�/�/�/�/�/	?.?  ������[?u�%-?ir�ectories ?�?�?�?�?�?O#O�5OGOYOkO��@ :�\\BKUP_1�9-JUL-24�_10-36-50\\oO�O�O�O�O �O__1_C_U_g_&=p��H?j?�_��!�?�5�Qdefr_oo +o=oOoaoso�o�o�o��o~�Full ;Sy�pm B;�o �o0BTfx`����+7���!�_�_�u�$�_�5�Summary/S0�^�p������� ��ʏ܏� ��)/;/ H�Z�l�~�������Ɵ ؟���� ��_�S�e�'�9�S1%���į ֯�����0�B�T� f�}O�O�O����ҿ� ����,�>�P�b�t��3�E��Ϲ���net�work��AutoDHCPy� �� $�6�H�Z�l�~ߐߢ� ������������
�� .�@�R�d�v����@���
�Ϝ�����&�����/roboti �o[�m���������� ��������3EW i{�����������1[�y=-�?�statu �?�����// ,/>/P/b/!a�Qg/ �/�/�/�/�/�/�/? "?4?F?X?);�?��?u�}�cllb ��j?�?OO&O8OJO \OnO�O�O�O�O!�O �O�O_"_4_F_X_j_ |_�_�_�_�Z?�?��_o��}�gripper�?AoSoeo wo�o�o�o�o�o�o�o �O+=Oas� ��������_��_�_0�Z�x�����2 �����Ώ������(�:�L�^�y�Fu�ll Sy��m B��c�������П� ����*�<�N�`�{ϐa�C����� y��s�ettingsp ������/�A�S�e� w�������ѿ��� ��+�=�O�a�sυ� �ϩϻ���� �r|ԯ�/name�� S�e�w߉ߛ߭߿���������r�ROBOT�5�G�Y�k�}� ������������� |?����R�l�&!o��ToolNum/Fr?�UsAߧ��� ������%7I[r�1_��� ����'9K]��
!�;���;��n)q���Active��b�/#/ 5/G/Y/k/}/�/�/`
0xf�$�/�/�/ ??*?<?N?`?r?�?�?�?�:�������?����Macr}o��s/New/B 5oROdOvO�O�O�O�O��O�O�O_�0x0_/_A_S_e_w_�_ �_�_�_�_�_�_o�60'��?CoUo�,O+K/BOpen���o�o �o�o�o%7I _r����� ���!�3�E�W�n��:o��
K-moooClos������ 1�C�U�g�y�����\�ԟ���
��.� @�R�d�v�������k�"}����N��/�Set/B��D�V�h� z�������¿Կ���YYeAO*�<�N�`� rτϖϨϺ�������4߼ �!���+o��G�	��'�ethodߙ߽߫��� ������)�;�M�'�Direct �entry of� EOAT dataW�������� ����%�7�I�߼! �"�4ߖ�M$i�'��traightOffsetZ��� (:L^p����"�� ��� �%7I[m ��b��v����BM%������%%X� G/Y/k/}/�/�/�/�/p�/�/�/�.00 �/)?;?M?_?q?�?�?@�?�?�?�?�?Oů�� �AO//'+Y O�O�O�O�O�O�O_ _+_=_O_?s_�_�_ �_�_�_�_�_oo'o 9oKo
OO.O�oROdOvOtZVo�o% 7I[m��b_ �����!�3�E� W�i�{�����^opo�o�䏦o)�o��Rot_ation!�W�� G�Y�k�}�������ş ן韨��1�C�U� g�y���������ӯ� ����ȏڏ<����"�nP��������ѿ� ����+�=����s� �ϗϩϻ�������� �'�9�K�
��.���R�d�v�nRR���� �%�7�I�[�m��� P�b����������!� 3�E�W�i�{�����^ߐp߂����k"����t�p3Zdir/Tp3z��<N`r ��������� &8J\n�� ��������������C/�`+	��Me�asuremen�t/Straigh�o�/�/�/�/�/�/ ??'?9?�
o?�? �?�?�?�?�?�?�?O #O5OGO//*/�ON/�`//We�!Num_s/New�CsNO �O�O_#_5_G_Y_k_8}_�_N=0xc?�_ �_�_�_o o2oDoVo hozo�o�ob@aO�i�O�o��.�O�LTo;ol�CUse�oD Vhz������Q:1��+�=� O�a�s���������͏Hߏ�a
�owD�o�1��o�LPart *������şן��� ��1�C��2G�m� �������ǯٯ���@�!�3�E��rI#�䅿��(Y��Gs/G ���CJ����
��.� @�R�d�vψϚ�]?�� ��������*�<�N� `�r߄ߖ�YOkO}O�����)����Payl?oad1CmԿ:� L�^�p�������������EOAT? w/o p{��� !�3�E�W�i�{����� �������������o 7���x����� �����0B�10��j| �������/`/0/B/��?	A ���/��W�2'��/�/ ??(?:?L?^?p?�?t�?���ith� �?�?�?�?OO1OCO UOgOyO�O��\/�O��OP&�/�)Advanced�O4_F_ X_j_|_�_�_�_�_�_�_��0x]o$o 6oHoZolo~o�o�o�o�o�o�o�@�O�O	�3M%�O�!Mas�s/Center gq�o������ ���)�;���_�q� ��������ˏݏ�� �%�7�N/��|�>�/bsssB�ߟ� ��'�9�K�]�o��� @�R���ɯۯ���� #�5�G�Y�k�}���N��`�r�ԿF,���!GPcmr��X��6�H� Z�l�~ϐϢϴ����� ����� �2�D�V�h� zߌߞ߰������ߥ����ɿ+�����sY �ߊ����������� ��,�����b�t��� ������������ (:����A�S�e�sZ>�� &8J\n�?�Q� �����/"/4/ F/X/j/|/�/M_q�/��.���1��$� 3?E?W?i?{?�?�?�? �?�?��OO/OAO SOeOwO�O�O�O�O�O �O�/�/�/(_�/�/?rtx�_�_�_�_�_ �_�_oo)o�?�?_o qo�o�o�o�o�o�o�o %7�O__|>_P_b_rt��� ��#�5�G�Y�k�}� <oNo��ŏ׏���� �1�C�U�g�y���J�\nП��|TCPVerify/
�?Method��.� @�R�d�v����������Я��Direct Entry߯ �"�4�F�X�j�|��� ����Ŀֿ������ȿ�!Ϗz'��fy "?|ώϠϲ������� ����0ߛ�T�f�x� �ߜ߮���������� �,ϻ�q�3�E�W�fyv_������� �*�<�N�`�r���C� ����������& 8J\n�?�m�c�0�����fy�$ 6HZl~��� �����/ /2/D/ V/h/z/�/�/�/�/�/����?���fyW�/y?�?�?�?�? �?�?�?	OO-O�QO cOuO�O�O�O�O�O�O �O__)_�/�/?n_0?B?T?yP2_�_�_ �_oo'o9oKo]ooo �o@O�o�o�o�o�o�o #5GYk}<_�N_`_��_�_�_yR �!�3�E�W�i�{��� ����ÏՏ�o���� /�A�S�e�w����������џ�����}*���fyMean ڟx���������ү�0����َ*?�+� X�j�|�������Ŀֿ �����ݟ�M���m��z)=�O�a�ax .���������%�7� I�[�m�,�>��ߵ��� �������!�3�E�W�i�{�:�|�^����{"��ϣ�Introductiof��)� ;�M�_�q��������� �������� 2 DVhz������������r�#��file2/�cyclepow��done�m �������/ !/��E/W/i/{/�/�/ �/�/�/�/�/??,;A��G?q?�r,���crsgdeta�il��Selec�tCategor?y/list,?�? �?�? OO$O6OHOZO�lOیAlloc��0d by KAREL{O�O�O�O�O �O__0_B_T_f_x_
�����Qw?Y?�_��|/�?��_for�ce/F�QLimit1�?o.o@oRo�dovo�o�o�o�oَ--- �O�o
 .@Rdv��� ���T�R�_�_��_�_�_`2op����� ����ʏ܏� ���o �o#�Z�l�~������� Ɵ؟���� ��!�`�e�'�9�K�t3_� į֯�����0�B� T�f�%�7�w�����ҿ �����,�>�P�b� t�3�u�W���{�����t4���*�<�N�`� r߄ߖߨߺ�y����� ��&�8�J�\�n�� ��������ϫ���+6����payl�oad�4PK�No?/check��x� ����������������  �OEWi {�������������^ �7�1�C�ldchg/�P�Enable?Signal�� ���/"/4/F/X/ j/�O;�/�/�/�/�/ �/??0?B?T?f?%
�Pb�PoQ�?!�����spdlmt�/S�2Clamp ��O-O?OQOcOuO �O�O�O�O���Њ/ �O__%_7_I_[_m_ _�_�_�_�_��?�?�o�78�?�5tat�us/SGbSafety�1
Oqo�o �o�o�o�o�o�o ~/�OI[m�� �������_�_��_<�f�(o:oLol2 `oŏ׏�����1� C�U�g�&8������ ӟ���	��-�?�Q� c�"�4�F�����|�����l3���+�=�O� a�s���������z��� ���'�9�K�]�o� �ϓϥϷ�v�������0�Я���l4�m� ߑߣߵ�����������E-�@ۿ@�R� d�v��������� ����������]��1�C߱5\������� ��	-?Qcο 4������ );M_�0�B�Ȍ��19}���usDigitalYo /!/3/E/W/i/{/�/ �/�/p��/�/?? /?A?S?e?w?�?�?�?�?~c���?O� ����iO{O�O�O�O �O�O�O�O_�/�/A_ S_e_w_�_�_�_�_�_ �_�_o�?�?�?4o^o  O2ODO��o�o�o�o '9K]_._ �������� #�5�G�Y�o*o<oNo ��ro�o�oW���1� C�U�g�y�������n ����	��-�?�Q� c�u���������|��� ���ď֏菩�_�q� ��������˿ݿ�� ��ҟ7�I�[�m�ϑ� �ϵ����������ί���T��(�:��6 U�����������&� 8�J�\��-ϒ��� ���������"�4�F��X��)�;߅���q�)�u߇�atsts/}A��Checkf� '9K]o����d�DISABLE ��� ,>Pbt����k�d�����/�+����TimeLm��X/j/|/�/ �/�/�/�/�/�/�� ?B?T?f?x?�?�?�? �?�?�?�?O�	/��MOg�5///InputA$�߲O�O�O�O��O__0_B_T_k�-- z�_�_�_�_ �_�_�_oo)o;oMo@_ov�0OBO�oj�0qO��OWarning �O%7I[m���f�x�s��) ����(�:�L�^�@p�������eo�pˁ��o�o�e�*�o�fr�sm��4�Enable��T�f�x����� ����ҟ���??� >�P�b�t��������� ί���O��I��g�3�+�PrgRun�o����̿޿� ��&�8�Jϵ�[� �Ϥ϶���������� "�4�F�X�ooY�;����cJ1m����Pause�����"�4�F� X�j�|���_�q��� ������0�B�T�f� x�������m�ߑ����eH%���c/Int�roduction��K]o��� ���������5 GYk}���� �����΁�����C/aL!'CompletB��/�/�/ �/�/�/??*?<?N? �?�?�?�?�?�? �?OO&O8OJO��/�-/wO�O�)i/�df/orce-F�AZO �O	__-_?_Q_c_u_ �_�_X?j?|?�_�_o o)o;oMo_oqo�o�o@�ofO�O�O�o^�/�O��J�BLimit1/var1�oQc u������� �_�_)�;�M�_�q��� ������ˏݏ���o@�o�oF�,{2; ����ğ֟����� 0�B���S������� ��ү�����,�>� P��Q�3���W�i�{�t3������*�<� N�`�rτϖ�U�g��� ������&�8�J�\� n߀ߒߤ�c�����������Ͽt4�H�Z� l�~���������� �ϻ���2�D�V�h�z� ���������������ߐ����=��.��JEscap4s7���� �����0 B��x���� ���//,/>/P/ !3�/�+a�JSummary�O �/�/?"?4?F?X?j? |?�?�?_q�?�?�? OO0OBOTOfOxO�O@�O[/�//�O��(�/�Comp�/=_O_ a_s_�_�_�_�_�_�_ �_�?�?'o9oKo]ooo �o�o�o�o�o�o�o�Op�O�O�OD��-	_��payload/IntroPws �o������� �+�=��_os����� ����͏ߏ���'��9�K�
.���5�]o|Select�tNo7����(� :�L�^�p�����S�e� ʯܯ� ��$�6�H� Z�l�~���O�a�s������3��o|�tWeigh��H�Z�l� ~ϐϢϴ������ϩ� �� �2�D�V�h�zߌ� �߰������ߥ���ɿ��=�[0��yqXYZ3ϕ������� ����%�7����m� ��������������� !3E��(��Py4Y�k�yqInertia���� #5GYk}�N� `�����//1/ C/U/g/y/�/�/\nȀ�/Tu/�Ýummary�:?L?^? p?�?�?�?�?�?�?�? ��$O6OHOZOlO~O �O�O�O�O�O�O�/�/��//_M|,?o|Comp)?�_�_�_�_�_��_�_	oo-o?nb �?Ovo�o�o�o�o�o��o�o*<�1mers__'_�KV�+U_gUldchg/IntroP�r A��	��-�?�Q��c�u����8gToo Uogȍޏ����&��8�J�\�n�����  timeWi{ݟ�KV1��{�sLimitX�:�L�^�p����������ʯܯ�7  ������ �2�D�V�h� z�������¿Կ��O��ɟ+�����#�Y )��Ϡϲ��������� ��0��?�f�xߊ� �߮����������� ,�>����!σ�E�W�i�tZ}������� *�<�N�`�r���C�U� ��������&8 J\n��Q�c�u���IX6���!�Rot����;M_q� ���������/ %/7/I/[/m//�/�/ �/�/�/���?0?�NS-��{Summary��?�?�?�? �?�?�?OO'O9O� 
/oO�O�O�O�O�O�O �O�O_#_5_�/"??�z_�}*M?�{Compt?�_�_�_oo0o BoTofoxo�oIO[O�o �o�o�o,>P bt�E_W_i_����+�_�Tspdl�mt/IntroS��1�C�U�g�y� ��������ӏ�o�o	� �-�?�Q�c�u����� ����ϟ០��&��Y2���Value/rw+���� ����Я�����*� ���`�r��������� ̿޿���&�8����	��}ϗV7I�[�m�tClampEn7abls�fl�_�� ����,�>�P�b�t� ��E�W���������� �(�:�L�^�p��A�0S�e������5�ϯ��mtMaxSpeedt�0�B�T�f�x� �����������ߣ� ,>Pbt�� ���������% C?��c�n3�}�� �����//1/ ��g/y/�/�/�/�/ �/�/�/	??-?� r?�_F��Ql�? �?�?OO(O:OLO^OpO�O4C/U/�O�O �O�O__&_8_J_\_ n_�_??m?c?�_��?>�tatus�b �_)o;oMo_oqo�o�o �o�o�o6/�O% 7I[m��� ���_�_�_�8�_ feoz������� ԏ���
��.��o�o d�v���������П� ����*��+��o� �?C�i�2i�˯ݯ� ��%�7�I�[�m�� >�P���ǿٿ���� !�3�E�W�i�{�:�L��^��ς�)���4atstdAц�#�5� G�Y�k�}ߏߡ߳��� ��������1�C�U� g�y��������� �϶���_����e� t��������������� (����^p� ������ @$����i��(=� �ʹ1c�����/ /1/C/U/g/y/8J �/�/�/�/�/	??-? ??Q?c?u?4FXz8�?��L�rsm� @ �?O1OCOUOgOyO�O �O�O�O�/�/�/	__ -_?_Q_c_u_�_�_�_ �_�_�?�?�?o.��? �7\�Oro�o�o�o�o �o�o�o&�O�O \n������ ���"��_#oog� �;o�8�aoÏՏ� ����/�A�S�e�w� 6H����џ���� �+�=�O�a�s�2�D��V���z�'��O�/S�electC��gory~��+�=�O��a�s���������Ϳ ��������,�>� P�b�tφϘϪϼ��Ϡ��˯����<&�n�etwork�s�ettingsp2/ipadd�� l�~ߐߢߴ����������� 
10.7� ?�D�V�h�z�� �����������
�� ��	���a��>ᯣ &����������� 0BTfѿw�� ����,>Pbt��;�M�����2��guid�ed�NetDone|
//./@/R/ d/v/�/�/�/�/}�/ �/??*?<?N?`?r? �?�?�?�?�?����O��5���Port�?\OnO�O�O�O�O@�O�O�O�O_�GA� 1 (CD38A)_R_d_v_�_�_ �_�_�_�_�_oo��W ���O��?_o}�1O��curit��o�o�o�o �o1CUg���?��Low �(R-30<i>�i</i>B S L�@_��������1�C�U�g���o-+ca3d���ooQo�����os/methoZ���)�;�M��_�q���������'V �= n�Man?ual icß�� ��+�=�O�a�s���p������̗1073dA��1Ï���%�ُ>�bummar�oZ� l�~�������ƿؿ� ���͖)��/>�P�b� tφϘϪϼ����������  eatu ;a�?�;�e�'���TesJO�������� ����,�>�P�b�#� en-ϒ����� �������"�4�F�X�~j�  tech'PA3�Eߏ���� ���s�tp1m� *<N`r����ђope���� 
.@Rdv�����  ageA(/ߕ���	/{f��>�Intro�U/ g/y/�/�/�/�/�/�/x�/	?'V800)� :?L?^?p?�?�?�?�?��?�?�? OO  penV���]O{f�%)/��/name O�O�O�O�O�O__�1_C_U_g^g() �ROBOTg_ �_�_�_�_�_�_oo`%o7oIo[oȞ u��gOIO�oq�&}O�Lipad�+=�Oas���l�i�gh�192.�168.150.2����'�9�K��]�o���������u�� o�o�o�w�'�o�Lsub5���]�o��� ������ɟ۟�����59-1�255.'�0�E�W�i� {�������ïկ����z�m',ӏ����Y��-��Drouter���ÿտ������/�A�S�c�0);
�{���Ϫϼ��� ������(�:�L�^�w�ady'�9�K���r&$y��Lmace� ��&�8�J�\�n�������72, ��00:e��4:�7d:bc:db ������'�9�K�]��o��������� {
  {ߍߟ�o����B2E�Rdv��������Addr %�2DVh z������� 
/y`��������U/ );���/�/�/�/�/�??%?7?I?[?@Q?uer�  �x/ �?�?�?�?�?�? OO�$O6OHOZOoSn=mi#/5/G/�O��}/; ���O__1_C_U_g_ y_�_�_�_xa�P���O �_�_o"o4oFoXojo�|o�o�o�o  ><�imwO�O�O�ok&!��Efile/ba�ckup��Summary�oOas ��������m�4��` �2�D�V� h�z�������ԏ���
�m��o�o+�U���B"/uprogress�����ȟ ڟ����"�4�F�X��R0���������ʯ ܯ� ��$�6�H�Z�_  
[ ��#��5�����B#�O��N�etTest/ipadd]����� /�A�S�e�wωϛϭ�� s)[]�1x82������	��-� ?�Q�c�u߇ߙ߫��V �o������k&&ſ׹linkstaG O�a�s�������������AR-2��	Connected "�'�9�K�]� o��������������� ��������D�v!�3�url��� ���/AS�g0WARN�h?ttp://�χ ������//)/;/M/�[3-?�/�m��Y/�/�/ ??/?A?S?e?w?�?<�?�<" DAq��? �?�?OO,O>OPObO�tO�O�O�O�P000 s��/�/�O�,q�����6�OR_d_v_�_�_��_�_�_�_�_�0 ?" �31�Ao .o@oRodovo�o�o�o �o�o�o�oq/�O!K__1\7�� ��� ��$�6�H���12:0�26@_~�������Ə؏ ���� �2�D��'9��]o�s8 U�����0�B�T�f��x�������l?���	SYSUIF�.VA A DG� EATCH.VR�������/�A� S�e�w�����Z�l�~� �����?!�3�E�W� i�{ύϟϱ��������� �\���#�5� G�Y�k�}ߏߡ߳���h������ �@0ְ ��տ�I��p��� ��������� ��$�x6�H�[�IS ic� v����������������*<N  vis=�%�7�[� ����,>�Pbt��[�id="���� // $/6/H/Z/l/~/�/�/?  /celgy ��/�?&?8?J?\? n?�?�?�?�?�?�?�?[�dius?O0O BOTOfOxO�O�O�O�Op�O�O�O� dir�/ �/�/A_?h_z_�_�_ �_�_�_�_�_
oo.o@o��loc__ro�o �o�o�o�o�o�o�&8J  FAN _!_3_�W_�� ����(�:�L�^�pp������.00� Ə؏���� �2�D� V�h�z������qe�w�����$FM�R2_GRP 1���� ��C4  B]��	 �1��C�.�F@ Y�@��.�G�  ��Fg�fC�8R��q�?�  ����.��6�X�Ѣ�87�5t��5����5`+�q�A�  ���BH�o�%�O@S331���-�S�d�.�@.�z�p�d� ����ֿ������	� B�-�?�x�cϜ���_CFG ���TC�������
߬�N�O �E�169511�R�M_CHKTYP  ��������ROMY�_MI�N_��������J�X�SSB�Ì�� �/��������߰�T�P_DEF_OW�  �����I�RCOM^���$�GENOVRD_�DO����=�TH����� dZ�dC�_�ENB/� C�RWAVC������� �Q�H!���ТI��P�I\ٳI.��}������}�ȁ�r�w��E� ���OU���� ��A��A�<ڒ����?�������>��C�  %�P�'9B��#pD����ߤ�SMT����� ��Ч��$�HOSTC��1�������� 	��������e$Ugy� ��C����/��	anonymous/G/Y/k/}/ �/������//1 �$?6?H?Z?�~?�? �?�?�?�//-/O O 2ODOVO�/�/�/�/�O �??�O�O
__._q? R_d_v_�_�_�O�?O �_�_oo*omOO�O �O�_�o�O�o�o�o�o E_&8J\n�o �_�_�����Ao Soeowoyj��o���� ��ď֏����0� S�A��x��������� ҟ�'�9��M�>��� b�t�����ۏ��ί� ��'�(�k�L�^�p������ן����18736��"�D�%� 7�I�[�mϰ��ϣϵ� ������.�@�!�3�E�pW�i߬���SM���ӷ5޿������� ��+�=��a�s�� �������������'�9��
�ENT �1��	�  P�!ros pc�E�����!1�92.168.1�50.10��  !������������& ��Jn1�U� �����4� X-�Q�u� ����0/�T// x/;/�/_/�/�/�/�/ �/?�/>??b?%?�? �?[?�??�?�?O�?�(O�?�?^O!AQU�ICC��=O!���2�OqG1�O�O!
1���B �@�OrF�O�OOOP_s@ROUTERR_._�K�O B?PCJOG�_}_�!  ��^CA�MPRT�_�_!���_�YRTk_o/o��o !Soft�ware Ope�rator Pawnelmo!�G�0 3�oT�NAM�E !c�!R?OBCONT_N��S_CFG 1��c� ��Auto-sta�rtedŴFTP �yq�߹��� �����Y�4�F� X�j��{�!���ď֏ ������RdvW� ���n�����ß՟�� ����/�A�d��w� ��������ѯz߼�η ��R�C���g�y��� ����r�ӿ���	�,� ƿ��Q�c�uχϙϫ� � ����&��Z�;� M�_�q�4�.ߧ߹��� �� ���%�7�I�[� m������������ ���!�3�E��i�{� ��������V����� /A������ �������� =Oas��*� ���//Xj| ���/��/�/�/�/ �/�?#?5?G?Y?|/ �/�?�?�?�?�?�?,/ >/P/Od?UO�/yO�O �O�O�O�?�O�O	__ >O?_�Oc_u_�_�_�_�3RI/&_ERR� �z�_�VPDUSIZ  3P�^j@��T>�UO�LL ��_.@ � �I��` 6���UWRD ?�@u-A�  guest3V�ro�o�o�o�o�o.tS�CD_GROUP� 3�@| Dq�"IIFT~$PA�~OMP~ �~_SH~ED �~$C~COM��PTTP_AUT�H 1�.k <�!iPenda�n�g�~zF�!K?AREL:*���}KC�#�5���VISION SET�`��j��������
���@���)�K�M�_�\q�tCTR*`�.mB`Ζ3Q�
n��FFF�9E3��+DFR�S:DEFAUL�T�FANU�C Web Server0ZߐΓ�t Zold��g�y�����������TWR_CON�FIG �u��Q���QI�DL_CPU_P5C�3QB�.@3�� >ɰ��MI�N$�	q >��~�GNR_IO�Q�b3P4h�HMI_EDIT �{�
 ($for�lead	�0Z$�cu.� h���?straig̿���regi  n�e����labelϵ�if��E��?jump iD�޽�kakujiku��ϸ�	undef`�������ݑ($�� B�4q1�j�Uߎ�y߲� �����������0��T�?�x�c����2�ROS2,14�91296301�  069��/[����NPT_SI�M_DOi�s�N�STAL_SCR�Ni� � �TPM?ODNTOL6��L�RTY�3�$���.�pENB6�	s�OLNK 1�.k�p�������� |2��MASTEh����˒��SLAV�E �.kH D���SRAMCAC�HEPb�qO_C3FG��	UO���~�CMT_OP�8k�2j�YCL��
�_ASG 1����Q
 4Wi {��������////A/<*NU�Mc2i
�IP���RTRY_CqN�2�_UP� a����U �� �#�����̔�)��P0�?�.k ����F?X?j?|?�?�? ;�5?�?�?�? OO$O �?HOZOlO~O�O�O1O �O�O�O�O_ _�O�O V_h_z_�_�_�_?_�_ �_�_
oo.o�_Rodo vo�o�o�o;oMo�o�o *<�o`r� ���I���� &�8���n������� ��ȏW�����"�4� F�Տj�|�������ğ S�e�����0�B�T� �x���������үa� ����,�>�P�߯� ��������ο�o�� �(�:�L�^��ϔ� �ϸ�����k�}��$� 6�H�Z�l��ϐߢߴ� ������y�� �2�D� V�h���	������� ������.�@�R�d� v�������������� ����*<N`r� ������ &8J\n�! �����/�4/�F/X/j/|/�/(3TOIMER�#�!,�%��"_MEMBER�S 2��%��  $#5�"���),�'�/9� R�CA_ACC 3���%�!   �X�T�iT��"6�]2  7� 
 Q6��O 5i�a?S6!Y6��834BUF001� 3�@;= M��u0  u0MU��4��4��3N�0*�2 �4@�4`�4�4UN�4N�4N�4O�4UO�4ODODP�4�P�4PDPKE�4P��4P�4P�4Q�4Q��4QDQDQ�4Q��4Q�4Q�4R�4R��4RDRDR�4R��4R�4R�4S�4S��4SDSDS�4S��4S�4S�4T�4T��4TDTDT�4T��4T�LT�` `� L�4M�4M�4MDMD�92�?�?�? �?OO*O<ONO`OrO �O�O�O�O�O�O�O_�_&_8_J_\_n]M@'��Q�Q�Q�Q�_�_2�]3�_�U  �S�p�R�p�R  �S�b �b�b��t#c��t3c  ;cB��Kc B��[cb��kcb�]�`�t�cb��t�c  �c ����c����c���t �c���t�c���c� ��c��ts��ts "��+s"��;s"��t Ks"��t[s�p�ks�p �rS�p�t�S�s!�s �p��s�p��s�"61�CFG 3�@;� 4�!�% <� �	��"34HIuS�2�@; �Q1� 2024-0�7-19& %!;�$`�!	�E \�(l��r`�8\��@l�H\�Pl�T�����ůׯ���*X�`C���S�	�H�PZ�l�~�#h\�pl�Qx\��1��\��l�U�\��l��\��l��\���Q`�X� C��1R�	�c�u�`��r	�����X\���	�!f����`����$Ěϸ�Ͼ���}C�6 ��s���O�a�	��� `���x�	�����ӿ�}]����5O���+� =�+�a�O�a���o�	�@w߉����	����� ����������	��� �ߟ���@�.�@�t�b��Џ�	�s�����3 ���ܼ�����:��� L���[�	�?�u��� �P-�?�����	������ :M0���  � �2�hz�|���&  A�� i�W�����{����|�� 9 c�&�  d�P	�ds��">�'  C�ϕ� �/�/����8/J/�n/ ����[�����ߵ� |"?X/F?�!�|?�� �?i�{���?���O ��f?TO�xOS�e� ?���O�O,O_,_>_ b_�O=�pRd�J!���b @�b�P�b 40�b�p�b�P�b�P�b � �b���b� �b�o  2D2DV�� ����b��b��b �0�bLP�bTP�b�@�b �@�b�0�b �b �b  �b/�o�o�o�o�o c�`� `�s���x�  �o���/?^�p��� ����<�����)�};��?0�B�T�f�x� ��������ҟ�bq�O ��0�B�T�f�x��� ����,�bq�_���� �0�B�T�f�x�������CI_CFG �3�xk H
�Cycle Ti�me�Bus}y�Idl��^��min����Up�ƺ�R�ead��Do�w����� ����C�ount��	Num ������]ݱz�CPROG����xe�`�L�/softpar�t/genlin�k?xpath=�/wizard/�file/bac�kup/step�s^curren�t=omenup�age,1631,�� ������|���4ձC SDT_ISOLC  xi�� U��|�$J�23_DSP_ENB  H�|ai�?INC �H��V�A�P?�0=�̟�<#�
U��:�o ������X���b�OB��Cr���B����(�G_GR�OUP 1�H�}�"< �^�P��t��?�n����Q���� �� 6HZl��� ��G_IN_AUT�O�D��i�POSR�E0�B�KANJI�_MASK��
K�ARELMON #�xkf߱y1J�\n����ӭ����(������ CL_L� NU�Mv��$KEYL?OGGING�@}`�!���LANGUAGE xe�P �DEF�AULT ^!faL�G��������9�P`�P����p'�R�t� 
���q��p�#� ;���
�!(UTg1:\��/ �/ ??'?>?K?]?o?�? �?�?�?�?�r(9
O���; N_DISP �����������?LOCTOLc@�q�Dz~�Q��yAGB�OOK �o-d �4���1�1�@�R�� �O�O�O__,^?]{#��QY-V	�E�Ip���+�_O��B_BU�FF 2�H� �_2���_�B(���_�� Coll�aborativ �Vo%nmodovo�o�o �o�o�o�o�o3*�<i`r�SDCS ��ٟ��N\�_�h�����'��tI�O 2��{ ��\���~��`�p��� ������ʏ܏�� �� $�8�H�Z�l����������ȟ؟����;�E_R_ITME�d� i�{�������ïկ� ����/�A�S�e�w����������ѿsG>�S�EV� 4M:�TYPF�X�9�K�]����RST/�uSC�RN_FL 2�
I�~Ч�������`��+�=�n�TP �E�(�mMNGNA�Mr��EP"$DUPS�_ACR�����D�IGI���U_�LOAD-�G �%j�%	DF_T�BIN���`�MA?XUALRM"��mP��
0���_�P���  �COQ0�C/@��M��o�%�A�q�N�P 2��K ؠ�	(������ �=�O�2�s�^���z� ����������'
 K6oRd��� ����#G* <}h����� ��///U/@/y/ d/�/�/�/�/�/�/�/ �/-??Q?<?u?�?j? �?�?�?�?�?O�?)O OMO_OBO�OnO�O�O �O�O�O_�O%_7__�[_F__(�DBGDEF �{��q����T_LDXDIS�A��i�9�MEMO�_AP��E ?j�
 �Q��	o o-o?oQocouo�o0��FRQ_CFG k�{��SA ���@��c��<�td%��l�o�o�`��{�{nT*?p=/Ar **:Jr�� =Ox�o��u��� ���� �l_{�I�� �:�p�^�t���,( �Ǐ�䵏�ُ��� '�L�3�p�W��������ʟ��� ��$�&�I�SC 1�j�0p �r_l�nT�_��m_���߯0�B�_MST�R ����SC/D 1��]�ׯQ� ӯu�`����������� �޿��;�&�_�J� oϕπϹϤ������ ��%��"�[�F��j� �ߎ��߲�������!� �E�0�i�T��x�� ����������/�� ?�e�P���t������� ��������+O: s^�������� 9$]�M�K�a���ao$�MLTARM�bu��g� ���P���PMETP�U�P
����N�DSP_ADCO�L��P.CMNT6/ %FN8 </>'FSTLI]/N'
� ���.��a��/�$%POSCFz~'G.PRPM;/��)ST 1��; 4�b#�
L1X L5\?j7H?j?l?~?�? �?�?�?�?�?,OO O bODOVO�OzO�O�O�A�!SING_CH�K  `/$MODA�c�J����YDEV 	>�Z	MC:wR�HSIZE�]
���UTASK %��Z%$123456789 �_�UWTRIG 1�� l�U�oo���_8o���VYPvQ��T�SEM_INF� 1�${`)�AT&FV0E�0=o�m)�aE0�V1&A3&B1�&D2&S0&C�1S0=�m)A#TZ�o�dH4�a(o\�hAd�G���� �o��o �o�o�oe������ ��r㏞��� �=� ��s�&�8�J���Ə ���(��ПڏK�� o�V�����X�ɯ|��� ����#�֟G�~�X�}� 0���\�ſ׿������ ��1�����yϋ�>� ����ώϘ�	���-� �Q�c�χ�:�L�^� p��ߔ���N�;��π_��p��|��rOoDONERŠ/�3S���   ����P�SN�ITOR� G ?�P[   	EOXEC1TX�2^�3^�4^�5^��P`�U7^�8^�9TY� ����]���i���u��� ���������������P��������2��2��U2��2��2��2U222*26�3��3��3i�QR�_GRP_SV �1Ɖk (�A@�H���-q=����>����?{�=���cXWSTR��ȉg!T�  �#��3T>A��"]�)EW�f x�E�Q�\��,����Q_DX�y^)#I_ON_DBP�]*3Q��3Pk+Xn%�w+�3PZ��!��N 3P/w/� ,X-ud1bU�/�/?�QPG_JOG �����
3P2  :�o�A=���?�!I?[? m?61>�?�?��;�?`�;�0|23P�1@�O8O&O8F  �Q3P�3STAT ��Z.1L_NAM�E !�U�@��!Defaul�t Person�ality (from FD)�!�QRMK_ENOgNLY�O�CR2�� 1��x����A; d�?_ _2_D_V_h_ z_�_�_�_�_�_�_�_ 
oo.o@oRodovo�� G1�o�o�o�o�o�op'9K �o r������� ��&�8�J�\�n��� ������ȏڏ���� "�4�F�X�j�|����� ��ğ֟�����0� B�T�f�x��������� ү�����,�>�P�b�t�����<a���� ҿ�����,�>�P��b�tχkA�a@.���3?������P�� ���"�4�F�X�j�|� �ߠ߲���������� ����B�T�f�x��� ������������,� >�P��1�������� ������(:L ^p���?u���� �  ����d �>�8F�?��0}�z�f  �����/�A�/#/�� (0m/4},���	`��/�/�/�!�1A�B�/? ?�?5 =@?9�**���"��C��3�  ��� (EW8C�  ä0��?��?��?O�?O:Oe	 >O%OzOeO�O�O�O�O�?�  �O�K�$�MRR_GRP '1�� QP(��"� � ��"P-P @D�#  @Q�E,Q?���A��@I�@U���O�  ;�	lXR	� �X � �P�R�Q ��, � �P�S� K�o���R��]K���K]�K	�.��Lv_�od�P@
�(baP0i�_�S��I�Xb�����T;gXb{Sў�]�3���b�1>�0�a�òN?v�?��=ڵ����?o0�o�bYQ�cT7�oUZ5�o } s��(p �  �  �8v�OV��U	'� � �trI� � � �L5�V:�����È=����u�R@��p�^2Q�BK2RD%��WyN� B�  'X�%aY`h�a`@e`h�mo#C�`���0C�`���m����"�_�_�XB� ���!��/=�q���Dz�O;��o_�pJ�o����R�����ഒА G4P��ŕ��zj1�K$  (�`?�ffW�����C � =�O��Q8��e�s�>L�p�`TQ�Z	(����P��ř�Q�U��R
���� x�Q;�e�m좢KZ;��=g;�4�<�<�ʏ�$��C��2S��<0?fff�?�p?&R��T@{=0d�?��p� ��"M�YT�O����ǿ 6��T'���� ��D� /�h�SόϞω���rh��F� ���ϭ�"� ��C߽��v�ߚ߅� �ߩ���������<� '�`�K��o�{��� o_��=��a�*�u�N�0`�r���#��"�7&%�A��A���=���(��"���JH9��A���i�����q�� �����0�-�D1ſ0���� �l�`P�8,ȴA;��^@��T@��^5@$�?��V��P�z������=#�
���?��
=�G}�pm�{=����,��C'���Bp�����6���C98R����@\)���(��5pmG��p�Gsb�F��}�G��tE�VD�K.����I�� F��W�E��E���D��;.����I��`E��G�]zE�vmD���, �/P�/�/�/�/�/#? ?G?2?W?}?h?�?�? �?�?�?�?O�?
OCO .OgORO�OvO�O�O�O �O�O	_�O-__Q_<_ u_`_r_�_�_�_�_�_ �_oo'oMo8oqo\o �o�o�o�o�o�o�o �o7"[Fj� ������!�� E�0�B�{�f�����Ï@���ҏ����(��34�]�ء���P��8�N��3~�qml�~�`��5Q����`���ğ֟������0���T�B�x�f���P�P������ӯ&�߯	�x��-������3� :�s�^�������Ϳ�� �ܿ� �9�$���0��cϙχ���Ϧ� ������� �6�$�Z�@H�~�lߎߴ��26���  B�R I ���CH"zm  @ Y�0�B�T�f�x���� H!���Т������l���?�� 

����Կ������
 �e�w� ���������������+=O����������U�$M�R_CABLE �2Ք� ��T������� ���� ������� Nt6H~�� ���/��/J/ p/2/D/z/�/�/�/�/ �/�/�/�/?F?l?.?� �*���?�?��?�?O#O5O��*XO** �O�M ו	�����*�h�?%�% 234567O8901�O�E �OH�O�A*��*��*��*�
�G��not sent� aJ�CW���TESTFECS�ALGR  eg���dZT3��A�lRà���*�o����_�_�_�_ 9U�D1:\main�tenances�.xml�_
o  �B��DEF�AULT��GR�P 2�yJ  �*���*�  ��%!1st cl�eaning o�f cont. �vPilatio�n 56�Bڦc �a�o��+A@���o`�o**�%�a�mech�`cal� check0  �js�tq{���o������?v�arollerRdv�k�l�~�𐏢���?qBas�ic quarterly�)�;��j,[�(�:�L�^�p�7ycMI��*�"8��!*���ǟ����� ��*�<���C�f������㟸�ʯܯ�� �?qOverghau�����>�C x*�H�O�����@|�������Ŀ*�$m� �Oۿ��k�@�R�d� vψ�׿�������� ��*�<�Nߝ�r��� ���Ϻ��������Q� ��8��'�߀��� ���������M�"�q� F�X�j�|������� ���7�0BT ��x��������� �i>��t ������// Se:/�^/p/�/�/ �/��//+/ ?O/$? 6?H?Z?l?�/�?�/�/ ?�?�?�?O O2O�? VO�?�?�?�O�O�O�O �O5O�O_kO_�Od_ v_�_�_�_�O�_�_1_ oU_*o<oNo`oro�_ �o�_�_�oo�o &8�o\�o�o��o �����M"�q �X��|�������ď ��7�I��m�B�T� f�x���ُ������ 3���,�>�P���t� ß՟矝�ί��� �e�:����������� ����ʿ��� �O�� s�H�Z�l�~ϐ�߿�� �����9�� �2�D� Vߥ�z����ϰ����� ����
��k�@�ߡ� v��ߚ�������W���	 X���-�?���B `�n������� ����������"4 FXj|���� ���0BT fx��������/n� Ў�?�  @��  L�G/Y/k/��3/�/�/ܼ/��*�/** F�@ h�j�  /?&?8?�/\?n?�?�?����]��/�? �?�?
O�?.O@OROdO �?�?"O�O�O�OO�O __*_pO�O�O6_�_ �_�_j_�_�_�_oH_ Z_�_Jo\ono�oBo�o��o�oo�on�����$MR_HIST� 2�f�"p� �
 \6�$ 23�45678901P2:t�o�"19/� ��Z�-���� ��E�W�i� �2��� ��Ïz�珞���ԏ A���e�w�.���R��� џ�������+��O���s���<�����pS�KCFMAP  ]f�%p�"�	q������ON?REL  ��"p�ڡpâEXCFE�NB�
أ��%�F�NC,��JOGO/VLIM�d"su��âKEY�x���_PAN������âRUNh�x��âSFSPDTY�PL��£SIGN|��T1MOTj���â_CE_G�RP 1�f� ڣ*r��/vσ�cϠ� Ċ��ς���߸�%� ��5�[���6�xߵ� l����������3�E� ,�i� �s�����z����������áQZ_EDIT	�ԧ���TCOM_CFG 1�Э/�|������ 
]�SI 	�M������������������W6�T_ARC�_)��W�T_M�N_MODE	�=�T�_SPLz:�UAP_CPL��;�NOCHECK� ?Ы �� "4FXj |��������//��NO_WA�IT_L�R�=�N�UM_RSPAC�EͯH�/�'�$?ODRDSP���7�OFFSET_�CARH���&DI�S�/�#S_A� A�RK	�S�OPEN_FILE� ����S���OPTION�_IO����T0M_�PRG %*%c$*�?�>03WO0[�M���p�5�i ����0��1	 ����3�f����� RG_D?SBL  wڡ�@/ORIEN�TTO���C���١A �"U� IM_D\7ע�� �V� LCT �@+�dt���I��d�i�C_PEX� �/�D�RAT� d7�|�D� UP �N
'p�`�\_n_T_�_��Y�$PALe���M��P_POS�_CH0_�QRA�M2F���x����C �@I%o7oIo[omoo �o�o�o�o�o�o�o !3EWi{���2o������ (�:�L�^����� ������Џ���� *�<�N�`�r������� ��̟ޟ���&�8� J�\�n���������ȯ گ����"�4�F�X� j�|�������Ŀֿ� ����0�B�T�f�x��ϜϞp<w������� ����0�B�T�f�x�|����kA�a�r��#�ߞy�P���ߞrP ���&�8�J�\�n�� ������������� "����X�j�|����� ����������0 BTf5�G���� ���,>P@bt������r	�!���KBd��/,-/N/\' ��F#�/��/�/|!�0�'�/�/�/�/?2A�'?9?�(��0h�?�<�r�%	`�/��?�?�?�1:�o��AOO,O>OG A��  UI�(@!@!ʞp"�pY$�~�C�  ����PPoFC�  ú@�/�O�/�O�O`___P_{%	T_�;_�_{_�_�_�_�_?�  �_k�$P�ARAM_GRO�UP 1�#0�(#K�� �2�� � �2~Fa @D�  Za�eFa?�pa�qC4�\cZa���_  ;��	lrb	 ��X  ��`�b�a �, � ��`�c~0�Hʪ��b����H���Hw�z/H��\�o�x",t~0B�  Bq�zaJyYs�3��rr�A>�@sq��ew�	�0B\�
��{�9�1K�^G"��rsa�jG�e�pE� }:���B�¨0�  �  �R��_p�u	'� � ���I� �  ��bEv=���8��ċr@ڏ�� ~La��;Lb^�?��wN@\�  'Dr�~0C�p���@C�p�������������B�o�oxB@
�A`�EM�2��1Dz�_�U��y�d�����r��Ƣ��΢?А 4PΒߥ"�5z�A?"����p??�ffm/�"��� �0W�i�q18�0���>LԀ�$naz(�0��Pĸߩ��a�e�b$���� x�}1;e�m¢K�Z;�=g;�4�<<��/�>��c�Lc��R@?f7ff?�?&l�t�@=0~�?����9Bg�sd�_�� ����PǦdA���:� %�^�I߂�mߦ߸ߣ� ���������6���� ��/��+������� ������2��V�A�z� e��������+��o�� W�{�D��hz���=��<�M6?�A��[�W<�'��d^I�;C�6�2-�%�3?���	��/� ��x`�@M$D1���J������!@�I�R,ȴA�;�^@��T@��^5@$�?�V+~0�z��ý��=#�
��� ?��
=��G�F-�{=����,��C'�?�Bp��� ���6��C98R����@\)��(��5F-�G�p�Gsb��F�}�G��t�E�VD�K�6>���I�� �F�W�E���E���D��;�6>���I��`�E�G�]z�E�vmD��� F/�?j/�?�?�?OO =O(OaOLOqO�O�O�O �O�O�O_�O'__$_ ]_H_�_l_�_�_�_�_ �_�_�_#ooGo2oko Vo�ozo�o�o�o�o�o �o1AgR� v������� -��Q�<�u�`����� ��Ϗ���ޏ��;� &�_�J�\����������ݟȟ���7�� (��!34�]9�����j�"�R�h��%3~��m����z��5Q8��įz���ޯ��!���
�
�J�@8�n�\�����P*�	Pľ�����@����#��G�2����� M�Tύ�xϝ��Ϯ��� �����/��S�>��`����}߳ߡ���� �������,��P�>�t�b������� 2<P���  B�lc��CH< zl� @ s8�J�\�n���������������6�#?�, 
$��#���� � ����
 � ������!�3EWi�*���������U�$P�ARAM_MEN�U ?
���  �DEFPULSE�@�	WAITT�MOUT�RC�V� SHE�LL_WRK.$�CUR_STYLv�,OPT"�N"/PTB7/1"C/R_DECSN� ��@܂/�/�/�/�/�/ �/??$?6?_?Z?l?�~?�?�SSREL?_ID  �ޱ���5USE_PR_OG %�%�?O�3CCR��2ޱ��G_HOST !�! D]OJoM_DA5 �
��Xe�.iU*HW2��=��7��lC��ETհ'O�C�@ORA�C�OK_TGIME��60E�?GDEBUG�0���3GINP_FLgMSK_GYTRV_�GWPGAtP 7\̼��[CHU_FXTY+PE����?�? o5o0oBoTo}oxo�o �o�o�o�o�o ,UPbt��� �����-�(�:��L�u�p�������IUW�ORD ?	�
? 	RSuPZ�/PNSX�$��sJON![�TE�@�COLXŹ�D�Z�WL�0 ��C���0Ed,QTRACECTL 1�G� ° �ݰ��ݱ����DT� Q�
�ِ��D � 	/���M �Y �U h��������,�I &�1ܱ�1��N���10�f�	�&�ݰ����6��� ��ʯܯ� ��$�6� H�Z�l�%�q������� ѿ����	��=�O� a�sυϗϩϻ�5��� ��%�7�I�[���o� aѭ���9����ݵ��� a��0�j�|�� �����~�H�Z����� 0�B�T�f�x������ ���������.�*< N`r����� ��&8J\ n������� �/"/4/F/X/j/|/ �/�/�/�/�/�/�/? ?0?B?T?f?x?�?�? �?�?�?�?�?OO,O >OPObOtO�O�O�O�O �O�O�O__(_:_L_ ^_p_�_�_�_�_�_�_ �_ oo$o6oHoRe& to�o�o�o�o�o�o�o (:L^p� ������ �� $�6�H�Z�l�~����� ��Ə؏���� �2� D�V�h�z������� ԟ���
��.�@�R� d�v���������Я� ����*�<�N�`�r� ��������̿޿�� �&�8�J�\�nπϒ� ho�����������"� 4�F�X�j�|ߎߠ߲� ����������0�B� T�f�x�������� ������,�>�P�b� t��������������� (:L^p� ������  $6HZl~�� �����/ /2/ D/V/h/z/�/�/�/�/��/�!�$PGTR�ACELEN  ��!  ���� ��&_U�P ����2!1)01"0�!_CFG �!5S3�!
"0�N4�N4h?s70s: � �s962DEF�SPD �A<��!0�� H_C�ONFIG �\!5	3 � � 5d�4�2 �!�1aP�4�1A� �� �IN90TRL ��A=a18�5 APEv�5��7�!1�N4�1�9LID:3��A=	|ILLB 1}��9 �E�B�0B4�Cs6 �H�G�OEu? �<< �!?� [-__%_G_u_[_}_ �_�_�_�_�_�_�_)oo1o_o|j�B�o�o �o�o_�o�o�o5~{IGRP 1��L��� @A!����4I��!A ��Cu�C�O_CjVF;|S0���4�1�y�y�1�0���@4_�A�~´���{B�/�����E�/�i�{�&�B34�����Ҏ��#Pj��׏�ӏ� F�1�j�U��y���u�x�ӟ  Dz� �R1��>��N�t�_� ���������˯�﯀�:�%�^�I�����)���
V7.10_beta1N4�0�@�*�@�) @�+A �2�?��
?ff�f>�����B�33A�yp0ͳB�(��A���AK��@kqxq 0˱ ˴̱�+�=�O�a�xqp����1l�ϥϱ�����R�fh����oB�!x�Z� t�z������%��p�$���4/rqBu�N� !5��� ����iA����lw� B�0B��ߦ��BH%��� ��r�G��Y1�W��x[�x�߁���������`0z�hB����������A�x����A�ff+��ia�DKNOW_M�  ~5I6�DSV7 ��:BS ,�������D����=�!�} A��*SYSTEM*� �V9.40341� {1/17/2�024 Ac�� h���@MSq_�T   � �$MAX_PYL�D�0$AXIS�INERTIA �  	$PSQ_�7�L� � ~�MOMENT��_� SC� � ��WT	INR�	  MN�.CL(PLD�_MODEDU_MMY11�0b�2j� MR� � $�_EN�B0$W}�^�ANGL]�@&}AA0�B���CC�DD�ST�_�,
$COM�P_SW�0�XOY_LO��Z%8� �� �� ����AYLOYA�7#_X=*Y=*UZ=*IJ+IX+If#�I�0DISP0��4� _RES�_G� | �5*SAV�� �)5�+6�%��&��&�2�#E�� UL0 �*}V�!  �@��$A�PMON�_QUE�!A@�$QCOU/!�Q�TH� HO�r0Hlj� IS~3UE]0=U�!�PO�@�!��$P[BU���OVERRU�N_TO�� O�DATA�!
@r�6C��CUR$�DEX�PROG�RA#� � 2N�E_NOD�5ITyPC�0INFO�!� �0�;/A��v31OI2B	 (0�SLEQ_NUMFC2@YP]qB�6�1�S_EDIT�!
3 �� K_�@kC$HIDE_� yU�G�HAUTO� �ECOPY�A�0�L�u$RMV_M�AN�@�Kv@�3PRcUT�t��NF�0UCH�G�21T�"�RGADJ�! �h� X_� I�1�$  ]V ]VW[XP�[XR[XSPEED�_MP�NEXT_�CYC�GSNS�_�3� $A�LGO_�0�NY�Q_FREQ�WqI�0wE�QSIZyC�1LAS�Q[Q#�P~kECREATE}3�0IFY�6NAM�]%,d_GSS�TATU� S�7MAILTIJ`p1wa�EV."�LASTxwa�!�TELEM�Q� ��ENAB<�`EASI�ap1 �� �bkA��f�;RO&0ATI@$��R�u1� rAB�1l`�0D_LV�a$vBAS~a$v�`�?sUPD_�0~`�$<qXwRMS_�TRs�� ts�S1P}3�aXt  �R�#� 	�b O2  b�	�`�wbr�w�rZ ��br�w6%�RARN_gDOU�3�IN���TPRE-P �aBGRIDA�3B�ARSjFP�cGROsTO� �! �1E_Hd!�Po�/�O�>�T � ��POR�3�����S�RVL`)����DIRECT_iҀ�Tu�3�4�5쉕6�7�8Ё�1F�Xq�1�0$VwALU?sGRO�2��d� �1F�U�C !�e��1��Na�0i�RAN��v�^a�R�@wAp1TOTAcL_{d
pԒPW�S�I7��REGEN���3Xex�3wE91���X0TRKsib�_!S�0K����cV[Qi8i�ukaGRE~c;��w1o2�2�@��V_H�X�DAX#k���S_�Y�Q��VSdAR�X 2 )RIG�_SEn3U����e_�0��C_c�$CM9P��DEV1 ݠ#�I�PZ���z+@F�HANC^1+� 
�g^byC���INTπ�QGF<�3!MASKZcVpOVR}3PO0;�t 8Ma�L�OVCbij:�AF9� 4f0H��jF%�c��PSLG��Q�r� �V� Z�ѐ|`S��d'�U��7I�}�V���`�eT$1O����CH���"!�l �r4 �*$�uA�J ��AC�cIL_Md��Vr�`�TQX0�3AR_pC'6�V�CݣP_��~`$�M;�V�1:�V1H�2W�2�H�3W�3H�4W�4 H��1i�r�1u���v�rIN��VIBhT��2�2�2�U3�3�4�4� � #Ԫ"��0�������������PLc`T�OR\0�p�Գ��B�RK��S�3�� ���bS� ^2d�� MC_F{0� �	e@����g�ǐMb+0Ig��� � �E"'�� KEEP__HNADD	�!K�$)pU�C*!L`k�o�
�� l�OQ1J��@�p�l�l�l�REM��k�{a��������U�Hdek�HPWD w K�SBM��~��COLLABZЗ�2�ő2bJ@IT��P��NO9!FCsAL�ēDON�R� ��$ ,0F�L�~a$SYN��yM����Q�U_P_DLY�!s�DELA� |a[bY�� ADX!$TA�BTP_R�4��QSKIP 	Ĩ��0O�u��r� P_�0�2 �0��  i%u%�$� $�$,�$9�$F��$9!q�RA�3� Xܠi���MB>��NFLIC�3���PU���7NO_�H� ���A��SWIuT2R�_PA @=G�q �!1b�UdpWJO�:#ߣg�NGRLT� �1{Q��K�M��<!�pT_�Ja&�rAP�W�EIGH�3J4CH�0a$ORu�a$��COO���b�a_&J����q�SA�!��#�(O�B�`�Y$)p!qz�Ji2�_1�EXJpT�S71#Aϑ71JPG��71AG� �RD�C��m ��@R����R!a��q���tRGEAD��`����FLG���0�(3�E9R��rSPC"C�Q�UM_70��2TH�2N2@�1 �4��o��R   D `��)-pW2_P�ECS[�|�q�PL10_Cbq!D�� !UP$K@мp�3�v�@���A�4�P�1���u�KA���CE`���r-s�  Fz�&@" P>,@DESIGbB�uVL1JI1WF�C	W;10��_DS���|�a;�POS11w�# l<�r�N�x�1#�/AT��"��U
8�RIND����}Q�SP��}Q`"�rHOM]E�R NOT2WR$]_o_�_�_�_�_`
PS3WR%�_�_�_oL"o4o �A�Q4WR&Woio{o�o�o�o�
PS5WR'�o�o�o
(.Fg6WR(Qc�u��� NU7WR)�����(�
@w8WR*K�]�o���L���� h0QPS >XQ+  ��PS���0C��K ��,� T,@]�ʖ]�IO���}�I���OK _�OP������1nCP�OWE��- �G�x U1�B�YP.�sؒ$DSB3�G#NA�B� C@���BMIc�/ ����)�1�0��P�$TP ɣ�෰W�AI�@>g KE � �3Y1�X��H�S�:��)ޡNEC-� 0� J��2�AL1Ʀ`AƢz�1t�OT�lS�1DLV�IC����W@QI߄SBN��% �PEA?��0�0���>20�ACC������H��5H�����1 `�]�U�F" [�UTOOL�\�M9UO�W2NC� R_��s�ANAD÷�b���2w2�BUFV���M� R�_VRS���IN �2@ӰH�0����(�_2 <�>����4�,�3Ǿ�A 3q0<�q�|�1 �@�S232c�3 ��y0ͅx�D�ICE�< �PE@�  I9T��OPB7 �oFLOW�TRa 0������CU��_��� UXT��4 T�ERFAC�İ�Uv���rSCH��4 t<��B�����!$FREEF�ROMW���GE:X I	�UPD"�iBf�1PT>�p%EX4��g�!�FA%�C��8 ��P�6�5+ &̈; A| �lى�0EX�IO#fрRY����_O��1P�����WR����D�1/�D��FRI,�z@�P����j���j�MYH�i�+�GTH_VTEY�1I�A��P$CPӰ~��UFINV_SP���H�RGI��f!ITI ��X�����G2��G1���@��<� �PRE_���<!DI"���#��t���ʐC> ��9�u�ALAR�0q$��Z� J���T�ҭ�$�� � 8% $�6�6 @n��0 ��Pd��"��$�A�� B���7�X ;"M��CT��H�@�0���Դ�G�3W�m��= �	D� ��Kq�� ϡ���A���� 2!6ʀ)�WP/�1;�*�U2-�2�3-�3;� �	-<��	I����L��!$VϠ��V��CV3����U�7�8w0#ֿ=�V2c��¹(�e�4�S�1E�0c���A���A����@�P!RQ0�pS����!ܒ��f�9 
P�1+� 740�� A8ʀ��:��@FR
@%�Sʑ: ؠR��!1�Bo�U��°X���S�ұL��NB�"T�H��I���@F�ER��4C�"IF_���&I-��#�� GA1(4�$9ĵ<67_JFE7PR�AIP��RVw; g $�A��  �BVALU�1Pj6zC�<Вx� 2; ��SCʒ=
  �$G�4A�2���4qT�@�#�3DSP�6�JOGLL���Y�P`0�5��!�3^@AXt�z�K}�_MIRAd!D9�MDBEAPc� E��&�1SYS�8A���1PGwFBRYKU��NC�0I�  �B.�B�2��qD{��3;@BSOR���3s�N�EDUMMY166i�נ����z�FC�_OVRi �HP�LDRCOIRW�NF�VF�!lV�0OVESFTZ� WSFpV2Q%C=���X����CHDLY�G=�OVT���0Wb��M���U@RO����A@_� �  @�d���VE_���OFeS��C�0Z�WD8Q��T4Q�Aق[E�@TRr��_�9�FDO[F�MB_CM��F`B�0BL�?�hb�+$�V$�o���3PRGig|HAMzC\`AЪe�R�o_M�`�9�x��PT$CA�09���>�T$HBKs��&qIO-�u��O�PPAz?q$yOt7u��e���RDVC_DB��q�!���p�R2Q"�u1�z�c�u3�v�PATIOF�0�QqU2��0x�CABY� ,�B�= �S��h�0�_
��&SUBCP	U��Z�S����Rc�d�t��S�p�d�Q$HW_C���䅇�A#� �$U�NIT�D����A�TTRI� ��Z�C'YCLC��A�rLC�FLTR_2_F�I4
��s��LP�K�4�SCT��F�_��F_��8���FqS���b��CHAF�� �y��b��x�RSD����������7p_T��hPRO�p@c��E#MP��@�CTf�wa��g����DI�О�$RAILP�/�MF�0LO�@���D7i�`��v��u�cPR�p%Sw�T�X�Ctq��=	�SFUNCR��RIN��s��AG�w���RA��t�R�Tp��D@	t��WAR53F�`BLq�ѤAʫƁͨƨDA갡��ѣʥLDd�P��4�d�!Q��3�TI��S��1� $/ RIYAHѽ�AFD�Pm�~��P��� �����MOIG�CfDF_�+��Sp���LM�cF�A��HRDY�ORG8�H��wQ'��>ҵMULSE+��#TS����JZJ6R�KWF[FAN_AL�MLV��R�WRNY�HARD�@s�����J�!�2Q����1�E)_�P��U��Rk��?TO_SBRvr����0�ʥ�vs���MPINF� ����)�n��REG.�NVq���ӚFDA��RdFL��R$M��%R�d�`� `�g�CM� uN� Y��NONI`��N�DEVY�j�s���� �I``�1>� �Y�$���$Z���2�1�0?o, �oCEG���3P�ѝ��t�E29pi����|EAXE�7wROB�:RED�6�W��A_]��CSYЯ@8�p�S��WRqI�P慀STR�5(���@*PE���0�C!3O �@����B���Qp��]��@�`OTO�9�0�PARY�3�0!��t�1AFI�@,C?$LINK���!J'�c_���Q��:�N�XYZw�Y��2!j�OFF�P&��N�B��B�0l�`���q̐p���FI)Р��w!R�Dl��4_JA�2(R3�;q����4��9!�TB���25C��kFDU��E�354�TURT�XZ�n���X��pFLm�P��� p�x���Ca 1>�0K�pM�$\3�S��S�%cORQɖ�1����84��@10ð�<p�#�1#�QOVEX�"M,�01��r��r ��q��o�p��o B5q�,����!Y9@� �r01jYv����L��1ERA �	8�!E�Pn0D�9$A�� ����Ē����AX�S�2�����(� �%���)��). �*e  �*�@�*3��*3�*!��*1���&���)���) ���)���)���)���) ���)��9��981,9x���~%DEBU}�$x�����1bJ�CAB�q8QRVp|� 
B�s!/E ��;G��;G.;Ge;G �A;G3�;G3;G!ኴp: �����LAB��qy��sGRO��4}��`B_ґ & ��͓�����FQU�� VAND� 8�.$ �qS�1!��]W �a�����qX��X�R�NT8d��S�PVELؑ���Q��X��͒��N�A�a��h�C��0%TRQL��Vvd���4�SERV9E�P��@ $��n�Q!1`POJ���_ĐT9�!	� b����A  #$Ub `�
Tch�2^`Bbg��2Aseb�~�_ C lT ���ERR���Ipp�P��aTOQ���L<��$���fĐG�3e%<�|"  TcR}E� D ,/a�we�`B�RAq �2C d8rfs��tj` E���$fג���"uOC|��`F  �k�COUNT�� �
��SFZN_wCFG]aG 4��%���T|#z��q�3�Q��aqp�q��H �,@Mz�+�!���oz��FAq����XX�5���a"G�4d̀X�Pz���H�ELAЭrI� 5��B_BASN|#RSR$�`�R�S<�L���1w��2�Ċ3Ċ4Ċ5Ċ6�Ċ7Ċ8w��RO0�Pq-�Q�NL��@�AB@c
���ACK�FINfpT_U�Up��	���T�_PUX,~�e�OUBcPà%����v����y&TPF?WD_KAR�a-�&�`RE?d�P#��EPQUE$�f YI �~���IU�C��O�p���P�O�SEM���G�EAȰA�STYfc�SO2�DDIo�����C�x'��_TM>9�MANRQ��O��ENDD$KEYSWITCH���Ǒ���HEI BE�ATM��PE(�L�E�bEQ P��UƓF�6�ǒS��DO_H�OM��Oz�W�EF9PR���rj��U��C�O���`qOV�_M��E��OCqM;�EA	 �;HK��J DL�&��pU�b�M�ᔒ�<FORC*�WA�R�1 !p��O}M� K @�4T���U��P'�1Ɣg��3�4Q���ESkpOא`��L$r�%�UNLO���d�b�ED��  ��S�@HDDN]aM� d`BLOB � � ��E�uN �<NЉ�y"��MS�UPGB��CAL�C_PLAN��1���AY���r���tOO � ��9 PI` $MѠ��5�B����Q-�Ml��C���ƹ�d��SC�eM�ЭQ�`@ aѹaQpt�Y|�Z|�EU�,��[��TaU��bе�rNP�X_AS�rP 0ί�ADD�p�q$�SIZ|!$VA�PuMULTIP�D����A��Q � $����F� ���М���C�`G�OFRIF��fpS���	�J�7�NF��ODBU� �PH���?f#CM��$@�1�C�t���.q��)`R g� ���bTE�\,3SGL�T5� &�p��C��S�TMT�5�PSE�G@�5�BWY�S�HOW=���BAN �TP����A�,0T�7ApTN�T>� S e �t	p���p��ALyI%b��OPENF��Q�q�WA��NEW_L�Õ���B��ز�q��RILN�_�BLK�P,P��- -EXp-SY�IPE��qJpF�TCz�B	�Ptx�Ʋ�� _BUFRQNW�� }�V+ �_G�rT 3$PaC�@gp+#�!FB��-P�SP�An����D� �rU�; ��aA00bT# �+'�+1�+;�+U5)6)7)8)9)A)��+�+ �A,��+� ++0�B51B���\1iU1v1�1�1�U1�1�1�1�U1�1�2(25U2B2O2\2iU2v2�2�2�@�`�(�Bp�(�2�U2�3(353BU3O3\3i3vU3�3�3�3�U3�3�3�3�U3�4(454BU4O4\4�94�9U4�94 I4I4�U4�4�4�4�U4�5(555BU5O5\5�95�9U5�95 I5I5�U5�5�5�5�U5�6(656BU6O6\6�96�9U6�96 I6I6�U6�6�6�Y6�U6�7(757BU7O7\7�97�9U7�97 I7I7�U7�7�7�Y7�i�7��rVD�_UP�DV��� 
��V��W x $TOR ������]�O�p'�t��tQ_�CURR��Z�AX(O�ҰZ�S�}C"���'�_� 1���YS�LO��X �  �Չ▣r���,��p%�<^�1�VALUh�y�H̖�q��FO�y L��ֿ�HI��I�$F�ILE_-�ꄽ�q$G��M�SAV�Y h�p�E_B�LCK��#�-�,�D_CPU<���<���������Y��k��R Z � �P: TO(���LA|SR�������RUN�Gŕ��ɑ���ʠ̕ꑷ�ꑬ�H`ด�����T2e�� ��[  $�JP���^�TPP_�EDI�$�S�PD,�\4�X�S|5����DCS���G�q] � $JPCQ�'�
7��S��C��C��$7MDL��$}�é3TC4�ŧUF�pĨ9SF�ĨCOB����T1��P����^� �����5������TABUI�_����_�� s]����^$���A���LB_AVAIY�� "���I�=`�p$SE�  ,1�DG_ɐN���
�pA* N�Ň�Q�!E� �����_}�.ʹ_��1�ELE�� ��SCRN Oa D��òB�T!ò�r��pN�Od�V�@�PRIO��t��VR��_MP��b \�pf�b 갤���M��D G� U4���6_�PS7��NѰ|�
�E̲��TBCD���c �̡C_BRK2_KMG��H�!�2+dW�e�B���Ď,�FTM��rf�2 �DC��C�б�`�L��x�TH}�u��Դ�ų�R�$��ERVEk���x������ BC_$� 2�c 	 �_AC��� eX -$�LENk��xӼ��RATI-�5$N�W��F1�ׄ2U�MO4���@��ERTIA��}��t���DE��8�LoACEM�wCCp�
#�V��X��������TCV����TRQ�#�����G�����J���p��a JH��������29�;������JK��VKk���x��������J0����JJv��JJ��AAL��P �� ��4 5��$�N1*�6 �����`t�
����CF���f `�pGROUP��v�f��N[�C�~� REQUIR��$DEBU����L�	��e��б ѫSGI�g��e�A�PPR��C�#�
u$=�NCLOr��S��)��
 �A;RA[�h �"�2����#��d9�1�GR��xL���y5�wN�OLDw��RTM!O+���hJ�@�P��������#���,�����7�8�=�}���J�i� ��5���T'x�b#PATH^'w!m#w!�:�s#T�h%�NT�e�Aj��mINF�UC��b�� CL�KUM�(YW���p �!Á���*��*��� �PAYLOA�J;2L�pR_A�75�L��C9?139O1xR_F2LSHR��|1LOD4�!}7�#�7�#ACRѠ�(�0�'�+4��H���$H�:��2FLEX�B!$�j Tr�MR 4���kDh4�Π:KeP� B7�ѲBJH�k l�W�i�����^��_FUN��W�E���j 	jA�l :�,���GT�/�ѱ�8�J�\�F1 QaUuWk�}������RE�������� )�;�M�_�|h�da��� ��c��h������Q��	T��zaX����X�� �W��Ju#h������  ��#,>Pb	���BJum � ����Q	ĐT��@k�U�0���a��J�vyAJE�CTR�ƊPTN)�\��HA_ND_VB BjA�OPoEn $�`F)2x���M��B|gCRo� $AdR���� H�& FA_.2hDU�qA�A�9Bz��H@��D�IB?I�XAGR�XAST�XB�XAN�DY�0x D�k�A0�s7Qs7�1@27���d;Pp�P� %%% %)%2%;#iB�oEp ��D\" ��Q��6�ASYIM�%=p�B�$o�P8�-�1�/_SHi�' �$�P�Ԉ�/??%?73J><�P:��o9.�T_VI��,�6>=�V_UNI��Q�ss{1J��j�j< nĥ5{ğƮ=k��9��?�?��+s�4 CK�E�CH�q�P |A��fTO/`PPp�V��B���
aR!PP��`eF�i�e�I�_�5!P�І��EѮ �RPROG_�NA�Q$a
$L�AST��cCAN�?P3�E�XYZ_SPA�U���)��}@�֑S"м���E�@��C;URd�FIR����?IO_TYP�cJ�GIND�G�.�X���E��@r@HR_TF�r͂����P���cO�����s �pr�J� j��  ��Pz���Pl�p �P��� t � �ME�Q� ���|�T��PTҰ]���p�t|@��"�=��1�TӰg+�DU�MMY1{q$P�S_�PRFNP�u$x���FLAw �N��%�$GLB_T�����3��@wLIF��u�R ��s�OW���d��V�OLw�.���_2�!g�2;!g���bا���+�TCyQ$�BAUDBQ��ST�BV�s�ARIT�Y<D_WAUAeI!	C��QOU�1�f�	TLANS���`SZ(�BUF_��@2`�J��CHK�@OCE�SUQr�JO�E����� ��UBYT�B�A�"^$:�m$����CY�B��S�CR�� v �.�E�P�P�R�PLUG������-����w L $PW3UP.�k�PWt��5L�Xk�EE�a��fIU����)�C_��PR����x� 8�0PIN5d�%6*7d�o���:"�yL d�����CH��,pu(OPEPNS� ��e����'��
e�2#�#-e�9e� Ae�O�"]�'3s�#�	�M1�	\7��M1�M1o��q�$��Q����z XX���pASTw����SBR��M21_�KХ`T$SV_E1R���5�3CL���2eA�POj�|�GL4��EW��{ 4 m$]�$a$�$W0C���ჯ�QRy�y�@UE|�{$��$GI���}$A {QTCI@��}�jGҦ�};ৱEsFNEsAR�P��$F�Ir�PT��� �J���RX� ~��$JOINT-q�p���AMSET�� E hGE�E�Q*�S1��UD*�����  ڊPU�Q?���LO?CK_FOL���oBGLV��GLdX�TE��XM��#QE�M w��R��OP�$US��@-p2|��IC�Q}yR�TP�Q�{�1CE�p|C�P �$KAR@aM��T�PDRA@�T�AV�ECLEj��DIUڮQ~�QHEVPTOcOL��+�#bVI,c;RE`IS3q?e�6�qn�CH	P9��*�ON#�<%#8`I�0� @$RAIL__BOXE-q��gROB�ЁR?��1?HOWWAR���a<u�jaROLM���e��qgd�b � :�ǀO�_F!�!��HTML5e�3�Q�܀1�E\a����N�e�TP:����BSLO�A�`��A� ��� t���U{|�f�u�OPr+POXq��I�ЂTN� 8b�b\a�ЮQ/p>��ORDEDTP9�LNp�@XT�pQ)G"���M� ��� D ��OB��j�TP�w��q�S���a |�YS�qADRk�|��!�>*� � ,π��'$A[Q��Y����BVWVA�� �� ��B��"R}T��$EDI��>��VSHWR�`�1�4�0�LAaH�Z��NBՃSHEADз����Ǳ��KE�a[�CP���JM�P	�L���RAC�E����pN�I��PS(�CHANN�E+`)��7TICK�,c_�M�z�/�H=N�1� @�pL�>�CP_GP�f���STY1�haLOB���B/������pp�
�Ь�%$~���=:�0S~�!$`�� ��N�M�PB��SQ�U�PޣLOO�+�T�ERC!���TS4�� r@��c�Dpr��a�#�F�IZ����L�t� ���4щ P�ʥ�_DO��X�X� S���AXI��b�Q.�&T�Њ��_��FREQ_`)�E!T*����\ AW��0!
�`H��ܰT�J�h�9��F z��SR_�1F��lj���p�RQ;s���$�0��B�ѳ�V�ѥ�/NOLDӹA]�A衷O���A��AV_@���ʿ��D�QD(�� <�J��C��C��)�C:���CY!Cn`w@��n`_"�������o�	tSS}C�� � hrpcDS����u`SPq�&�AT'���ˡ���X�d�ADDR��$T =IF�ӥP_'2CHL2!�I�0L1��TU�0I�� ���BCUO K��V
9RI��J�dX+�M�*�
�Z
G"VgqڡNF�� \��x������@��C[Ë�N�p�ڀv�2���TX{�EE�r���+ }PICNACy@I�Dv�8+�+�
Б T>��0 ����0�0����{#���䥀RR�A(���؏���+�UE4�� �������S	A)�RSM���U�pT��> �THRS_CC �@���#�>���+�CIR���}� 2�D�UE��� ���b��� GMTN_FL�g���0�q�A�@B�BL_l`W� F��S ����O=A��LE[���`����R7IGH�RD�4Q�OCKGR� T�p|WIDTH�3x��"�1FLAG����I�`EYpE��� d!@p�`̒� �aBACKʑ�b{��1u FO�q�L[ABձ?(u I*PMR$UR�a� T@�T MENH�� �"� T_�L2�؀R�OR�3rh���)Ob�F����GO0�U��,R]R�aLUqM,�&K�ERV�q�P�@[� � _�GE��AI��r&�LP~G�EQ��)�������V`�U5�6�7�8�@O������@
�te1�3� �SUS=RD� <��� 1UoB��oBFO��oBPRIg�mv`��} �TRIP�am��UN� 4��f@ �� 略a$��R(��0� ��H ��G ���T�`��M1�"O	Soa�&R.����#(a�A�O1C8N2���%�#U�A�?+?p9����#OFF~P*
О�A3O�0�Pќrp�4�4�rpGU#�P�1;r�3���7h�SUB�� �E/_EXE3�VG��#�WO�� �`0��'�WA��H Az�PG�V_DB*CHB@��H T0�������A�`��ORl`rERAU��sDT�IA�XAy_��4�� |���A�OWN�P`�$GSRC��H��D~P<�E��MPFIÔw�*�ESPơ��a�:e[}aWHb۫E����G� `b0B`���n/�COP�$�� _�@r�lQhqsU4BCTA&SAHb���~��b�� ���SHADOW�,c�Q?_UNSCAc�S�@�SDGDaa�E�GACfS���V�CͰCY3�� ��b"��$`EAR��/l-�t��Co^/eDRIV��5�C_V��Rd��a�D)$?MY_UBY($7d��3���.�a�ہ�h�Q�bP_�PÔ�bmLЫBM��$W�7DEYF�EX�p��wUMU#�X��"t�cUS���x _R_�@�m 
���A�G\�P�ACINg��RG �A[tqrw3qr63qrH�lQRE�_�1�28cqr
Х ��^P�Gw`P,�p� cR 0
Цc %��I�2�	kR�RE.sSW&ip_Ajq�0#s���O>!Q�Ac�*���E"��Uې� �1��c+HK���"B�B�0��'���s�EAy�}��@o@*�N0bMRC]V7�� �wO�Mo@C-�	���3�s��REF��܆Æ�� �hX��M ���Њ ��4�Æi�_�@�j����S w�cz�p�Abb}�� �𠈡�rN�Y!�el�O�U�3��r1�7c 3��u��2�#@J�๠���*�����l�K�ULW��+P3CO��fP�p�NT&SS��RR�^�5!^��L�c���c�����5!�VGR������ $�����O� ���BVL�O��$X������I��SY����QDO
x`EQ&#��c2��PIX�w31�SZ #��d^��d2�H��`h1�Q��B��SIb� l2��������}�f��  ^r~�a�Ipq۳Q���}�x�JvTZ�_AR�Y��o@REDU�Cs�FIT��P�RJвQ�l2LINE_XYSKI.s�M���5VIAF�� � @HDt�s �$JO ���?$Z_UPLy ��ZT���m�����_M�i�EP��#�)�� m�=�D�YD��l�)b��� 5*�P�A5 �CACHs���p8�@�P�CC��MI�SF���d�T��c֤�$H�Oo@�B!�COM	MMc��O���͗I`g�A�{єPVP�r ��Ѡ�s��ZUp�ذ����4AMP�F�AI��Go�2�A9DA�lRMREДa���GP�
p���S�YNBUFvVVR�TD��䠱OL�E_2D_q3��W.63PC_v`Us�yQG���ECCU�x�VEM�p��b�VIRCA�ś�ҟ�_DELA�s�A� �� �dAG��RqXYb��CqW�qs���F��1 �T`rIM�Y��;�@ W�GRA�BB1Y.s3�LE�R<pC���F_D�`��+&50������p�P(c��� �p��LASs���_;GEĥ� ����A$��TT���Aa,P�6"�uI{�r?�B?G_LEVEat`�PKtpA��A͗GID NO,Qq�qA O�$n�Я�"O�Sc�.�IN�T�LAŤ��R��Cױ`'#��D�!DE ��A:�P:�dp��  T�<��@�2��T  �-$5#�iJNQDq!�M1o T���ؑd@� $#AIT��"<��eSh�S9FaPƣ�  � 'k�^�pURrqSM�%��"�HADJ��u��ZD�� D���AL��`���޻�PERI��$�MSG_Q�$@���= 4B�d@�����!M������WN�`�D� � ����`�q �"`C��`0$�"�0�BJ4`s���Qpb@&6WN��C�XVR�C�|,�T_OVR'��ZABC_E���rg2���
 }�X!ACTVS��� � � $x�51q"CTIV屆��IOmb�3���QI�TcprDVP
Hpq�@�`,��A�0PS���B Z��B��8�p�1��LST�R��ر��1E_S�Q|<X!DCSCH�B� L�SD�5O�Pp���P����GNA���(@s��S@_FUN������ZI�%�L�	g$L����p_ZMPCFk5�"p�@6�A�aLNK�r�
�Ak�l4�� $��}�4CMCM���SC_Q.Q��P�1 $JLSFTD��RRcR\W �hU FWπքaR�WU9X~�5UXE)q�V ~�WU�UmU�Q�Q�Y�Q�WKPFTF?�RSd�e0�%��"<(�D�%"&aYM�D�� g� 8f�հIU)3�HEIGH\s�?( ��&����&`��� � �灅0�$B�t�uq�SH�IF��<(RV��F ���b\0C��GR<Q 0��Gr�aPS���YDx�CE0V��|M@߰PHEREч� , �ahwo�i��$��# 1 �����q���ДA p	 �pp3#�	��s�r�v��w�v��
]b�s7�@��q �q���� ���q�� k1�}T�uB�� 
 \�t���_���qN�BANFWD9 n�q�q���K ݰ1 1�u�߀p�4EO�AT w/o p�art_��� 	��r4��%�j�I�[� �����֟��ǟ�� ���!�3�E�W�i�{����ү��ɇ2Ԍ�q4>��  �<�寂ݰ3����1�ɇ4 N�`�r���ɇ5����ſ׿ɇ6����*ςɇ7G�Y�k�}�ɇ8`�ϬϾ���ɇMA���& ��  ���O�VLD  ��`���Ʉ�`�! ׋ r�HѼߎ�U@?و0N��
���!����UP�D��p�H�<�F�ɂ_�C� �! �p�'q��X���CHKf������rz�c�u�RSS����q������C@���y_GӀ��
 4���A�F�w� j��������������� =0B���"�2�d�M���� ������� #�F�>]b� ��}�������<��V 1�u��>�q�[�l��%0G_IN�0CҪqd���dO&MASS\/ �Zp'MN[/�#MO�N_QUEUE #�u������A*�N]�U��N�&�(��#END�!��)EaX@?�#@BE0��/�#�c�'�� eqR�AM %�*%�� /���"TASKhqN?��O A�/xrߵ?�0DATA�s]�;@�v2�u WOiO{O�O�OJO�O�O �O�O_�O/_A_S_e_^OINFO�s5M��$!_�_�_�_�_o o*o<oNo`oro�o�o �o�o�o�o�o&4�W�T	5L P	�1~~�DIT 
�?����4WERFL�-8B#��RGADJ7 uzA�Π�t�?��uc!�v�!�0}C��?���9z#&EA<@�R�V�%�T��xP�/A2Y�Ur	H� l#'yA"�>���Хw�t$Ć*Ӏ=/Ղ **:ނАя����u����С��qC�R=� �s��-�[�Q�c�ݟ ����ǟ��ϟI��� 3�)�;���_�q����� ��!�˯ݯ����� 7�I�w�m�������� �ٿ�e��!�O�E� W���{ύϻϱ���=� ����'��/ߩ�S�e� �߉ߛ��������� ��+�=�k�a�s��� ���������Y��� C�9�K���o������� ��1����#�@GY�}�:&	O (O:ŉqǃ�=�9���PR�EF ��
)$RIORI�TY�'�&��qMP�DSPk1�z�R/'U��'���vODUCT��1�zE169511��0���_TG�p�2yzn"HIBIT_DO-?�l$TOENT 1�u{ (!AF_INEY ?7?!tcp??=�!ud.?g>!icmV?]�n"kXY
�u|�Q�)� ��?�?��?O�5�?2OOVO =OOO�OsO�O�O�O�O �O
_�O._@_*m#
����RB��_�_<�>S�>�p��/��Hr_�_���j�u�A3�?,  � [q@0oBoTofo�u���V�Z�_�o�o�o�o�S�USENHANCE� a]_rAwkdx�_<#u  �j&��|& .v1�qPOR_T_NUMZ#��%�q_CAR�TREP� �<"S�KSTAY'�+SL�GS	0�;���SUnothingD%�7�I�Y���|���������pT?EMP })����m�_a_seiban���,� R�=�v�a��������� �͟ߟ��<�'�`� K���o�������ޯɯ ��&��J�5�G��� k�����ȿ���׿�� "��F�1�j�Uώ�y� �ϝϯ��������0� �T�?�dߊ�u߮ߙ���߽������,�  �$H ���sVE�RSI8 {'}� �disabl�eVp��SAVE �}*	267_0H705/����!,����h?� !	5�c"�g�^��S�e{���������������ro��_�  �1�;�� �}'I�l~�^�URGE�`B� �.�1WF� �!\$}b��&W0�D!�zWR�UP_DELAY� �}@&�_HOT %}%e"+�O�R_NORM�AL.�">�bS�EMIr��L!Q/SKIPJlw[x�/�@/R/d/'- Q�/�/�/�/�/�/? �/?7?I?[?!??m? �?�?�?�?�?�?�?!O 3OEOOiOWOyO�O�O �O�O�O�O__/_�O�?_e_S_�_�_�_]�RACFG ��l;���Q_PA�RAM�3�; Dzh@`�d�2Cp�;�@�Q�Cv�qBBH>�RBTIF�~�PCVTMOU�w��u��PDCR�J� ��3!?�ͦB?�"Bɳ@�5�?�8�;t�7'-�����Y�?����Sq*/�&.;e�m2r��KZ;�=g;�?4�<<�� 8p�} �� ������%�7��I�[�m��RDIO�_TYPE  �Qaw�EDPRO[T_�Q �B��0[a�EL`Ň�2�!Ջ �^qB� X`�*�^P�t�_� ����+�ɟ��{/� o_!�#�5�k�Y���}� ����ߟ�ie����� 1��U�C�e�g�y��� ѯֿ�������-�� Q�?�u�cϙϻ���߿ ���ύ���;�)�K� q�_ߕ߷ϼ��ϝ�w� ����7�%�[�I�� �ߦ��w���s����� ��!�W�E�{���� ����������� A/Q�����kcŇ?INT 2"1�=��aG;� ���;�[��f�0  4FcfWvx� �����//>/ ,/b/H/Z/�/�/�/�/ �/�/�/??:?(?^? p?V?�?�?�?�?�?�? �?O O6O$OFOlORO�O~O�O�^EFPO�S1 1#�� @ x�Y�c	 +__O_[X�O_A_�_ �_�_a_�_�_o�_o Do�_hoo�o'o�o�o ]ooo�o
�o.�oR �ovs�G�k ���*����r� ]���1���U�ޏy�ۏ ���8�ӏ\������� -�?�y�ڟş����"� ��F��C�|����;� į_���������B� -�f����%���I��� ��ϣ�,�ǿP�b� ���IϪϕ���i��� ��߱��L���p�� ��/߸���e�w߱�� ��6���Z���~��{� ��O���s���� �2� �����z�e���9��� ]���������@�� d����5G�� ��*�N�K ��C�g�/ ���J/5/n/	/�/ -/�/Q/�/�/�/?�/ 4?�/X?j???Q?�? �?�?q?�?�?O�?O TO�?xOO�O7O�O�O mOO�O__>_�Ob_ �O�_!_�_�_W_�_{_ o�_(o:o�_�_!o�o mo�oAo�oeo�o�o�o $�oH�ol�� =O�����2� �V��S���'���K� ԏo���
������R� =�v����5���Y��� �������<�ן`�r� ��Y�����ޯy�� ��&���#�\������ ��?�ȿڿu�����"� �F��j�ώ�)ϋ� ��_��σ�ߧ�0�B� ����)ߊ�u߮�I��� m��ߑ���,���P��� t����E�W���� �����:���^���[� ��/���S���w�  ������ZE~� =�a��� � D�hz'a� ���
/�./�+/ d/��/#/�/G/�/�/��$REFPOS�2 1$����1 @ x}/�/�/G?2?k? q/�?*?�?N?�?�?�? O�?1O�?UOgOOO NO�O�O�OnO�O�O_ �O_Q_�Ou__�_4_ �_�_j_|_�_oo;o �__o�_�oo�o�oTo �oxo�o%7�o�o j�>�b� ��!��E��i�� ����:�L����ҏ� ��/�ʏS��P���$� ��H�џl�������� �O�:�s����2��� V���񯌯���9�ԯ ]�o�
��V�����ۿ v�����#Ͼ� �Y��� }�ϡ�<�����rτ� ���
�C���g�ߋ� &߈���\��߀�	�� -�?�����&��r�� F���j������)��� M���q������B�T� ��������7��[ ��X�,�P�t ����WB{ �:�^��� /�A/�e/w//$/ ^/�/�/�/~/?�/+? �/(?a?�/�? ?�?D? �?�?z?�?�?'OOKO �?oO
O�O.O�O�OdO �O�O_�O5_G_�O�O ._�_z_�_N_�_r_�_ �_�_1o�_Uo�_yoo �o�oJo\o�o�o�o �o?�oc�o`�4 �X�|���� �_�J������B�ˏ f�ȏ���%���I�� m���,�f�ǟ��� �����3�Ο0�i�� ��(���L�կ篂��� ί/��S��w���� 6���ѿl�����ϴ� =�O����6ϗςϻ� V���z�ߞ� �9��� ]��ρ�ߥ߷�R�d� ������#��G���k� �h��<���`���� �������g�R��� &���J���n���	�� -��Q��u�"4�n��� �$R�EFPOS3 1�%��� @ x� ��dO���G �k�/�*/�N/ �r/�//1/k/�/�/ �/�/?�/8?�/5?n? 	?�?-?�?Q?�?�?�? �?�?4OOXO�?|OO �O;O�O�OqO�O�O_ �OB_T_�O_;_�_�_ �_[_�__o�_o>o �_bo�_�o!o�o�oWo io�o�o(�oL�o pm�A�e� ��$����l�W� ��+���O�؏s�Տ� ��2�͏V��z���'� 9�s�ԟ��������� @�۟=�v����5��� Y��������ۯ<�'� `��������C���޿ y�ϝ�&���J�\��� 	�CϤϏ���c��χ� ߫��F���j�ߎ� )߲���_�q߫���� 0���T���x��u�� I���m�����,��� ���t�_���3���W� ��{�����:��^ ����/A{��  �$�H�E~ �=�a��� ��D///h//�/'/ �/K/�/�/�/
?�/.? �/R?d?�/?K?�?�? �?k?�?�?O�?ONO �?rOO�O1O�O�OgO yO�O_�O8_�O\_�O �__}_�_Q_�_u_�_ �_"o4o�_�_o|ogo �o;o�o_o�o�o�o �oB�of��7 I�����,�� P��M���!���E�Ώ i��������L�7� p����/���S���� �����6�џZ�l�� �S�����دs�����  ����V��z���� 9�¿Կo������� @�ۿd�����#υϾ� Y���}�ߡ�*�<��� ��#߄�oߨ�C���g� �ߋ���&���J���n� 	���?�Q����������$REFP�OS4 1&����;� @ x������� l�������d������� #��G��k�� <N����1 �U�R�&�J �n�	/���Q/ </u//�/4/�/X/�/ �/�/?�/;?�/_?q? ??X?�?�?�?x?O �?%O�?"O[O�?OO �O>O�O�OtO�O�O!_ _E_�Oi__�_(_�_ �_^_�_�_o�_/oAo �_�_(o�oto�oHo�o lo�o�o�o+�oO�o s��DV�� ���9��]��Z� ��.���R�ۏv���� ������Y�D�}���� <�ş`�������� C�ޟg�y��&�`��� ��寀�	���-�ȯ*� c�����"���F�Ͽ� |���ȿ)��M��q� ϕ�0ϒ���f��ϊ� ߮�7�I�����0ߑ� |ߵ�P���t��ߘ��� 3���W���{���� L�^���������A� ��e� �b���6���Z� ��~����� a L� �D�h� �'�K�o� .h����/ �5/�2/k//�/*/ �/N/�/�/�/�/�/1? ?U?�/y??�?8?�? �?n?�?�?O�??OQO �?�?8O�O�O�OXO�O |O_�O_;_�O__�O �__�_�_T_f_�_o �_%o�_Io�_moojo �o>o�obo�o�o! �o�oiT�(� L�p���/�� S��w���$�6�p�я ���������=�؏:� s����2���V�ߟ� ����؟9�$�]����� ���@���ۯv����� #���G�Y����@��� ��ſ`�鿄�Ϩ�
� C�޿g�ϋ�&ϯ��π\�nϨ�	���-�:���$REFPOS5 1'���X�� @ x���� ߞ߉����� �߁�
���@���d� �߈�#���Y�k�� ���*���N���r�� o���C���g����� &����nY�- �Q�u��4 �X�|�);u ����/�B/� ?/x//�/7/�/[/�/ �/�/�/�/>?)?b?�/ �?!?�?E?�?�?{?O �?(O�?LO^O�?OEO �O�O�OeO�O�O_�O _H_�Ol__�_+_�_ �_a_s_�_o�_2o�_ Vo�_zoowo�oKo�o oo�o�o.�o�o va�5�Y�} ���<��`���� ��1�C�}�ޏɏ��� &���J��G������ ?�ȟc��������� F�1�j����)���M� ��诃����0�˯T� f���M�����ҿm� ����ϵ��P��t� Ϙ�3ϼ���i�{ϵ� ��:���^��ς�� ߸�S���w� ��$� 6������~�i��=� ��a������ ���D� ��h������9�K��� ����
��.��R�� O�#�G�k� ���N9r �1�U���/ �8/�\/n/	//U/ �/�/�/u/�/�/"?�/ ?X?�/|??�?;?�? �?q?�?�?O	OBO�? fOO�O%O�O�O[O�O O_�O,_>_�O�O%_ �_q_�_E_�_i_�_�_ �_(o�_Lo�_poo�o �oAoSo�o�o�o�o 6�oZ�oW�+� O�s����� V�A�z����9�]� ���������@�ۏd� v��#�]������}� ���*�ş'�`����� ���C�̯ޯy���ů�&��J�W��$RE�FPOS6 1(����u�? @ x�� =�����߿�Ϟ�'� ¿$�]�����ϥ�@� ����vψ���#��G� ��k�ߏ�*ߌ���`� �߄���1�C����� *��v��J���n��� ����-���Q���u�� ����F�X������� ��;��_��\�0 �T�x�� �[F�>� b���!/�E/� i/{//(/b/�/�/�/ �/?�//?�/,?e? ? �?$?�?H?�?�?~?�? �?+OOOO�?sOO�O 2O�O�OhO�O�O_�O 9_K_�O�O2_�_~_�_ R_�_v_�_�_�_5o�_ Yo�_}oo�o�oNo`o �o�o�o�oC�og d�8�\�� 	�����c�N��� "���F�Ϗj�̏��� )�ďM��q����0� j�˟������7� ҟ4�m����,���P� ٯ믆���ү3��W� �{����:���տp� ����ϸ�A�S�� � :ϛφϿ�Z���~�� ���=���a��υ� � �߻�V�hߢ����'� ��K���o�
�l��@� ��d�����#����� 
�k�V���*���N��� r�����1��U�� y�&8r��� ��?�<u �4�X���� �;/&/_/��//�/ B/�/�/x/?�/%?�/ I?[?�/?B?�?�?�? b?�?�?O�?OEO�? iOO�O(O�O�O^OpO �O_�O/_�OS_�Ow_ _t_�_H_�_l_�_�_ o+o�_�_oso^o�o 2o�oVo�ozo�o�o 9�o]�o��.@ z����#��G� �D�}����<�ŏ`� ��������C�.�g��t��$REFPO�S7 1)������ @ x� �Z�؟ß ��� ���D�ߟA�z� ���9�¯]������ ��߯@�+�d�����#� ��G����}�ϡ�*� ſN�`����GϨϓ� ��g��ϋ�߯��J� ��n�	ߒ�-߶���c� u߯����4���X��� |��y��M���q��� ���0������x�c� ��7���[������ ��>��b����3 E���(� L�I��A� e� /���H/3/ l//�/+/�/O/�/�/ �/?�/2?�/V?h?? ?O?�?�?�?o?�?�? O�?ORO�?vOO�O 5O�O�OkO}O�O__ <_�O`_�O�__�_�_ U_�_y_o�_&o8o�_ �_o�oko�o?o�oco �o�o�o"�oF�oj ��;M��� ��0��T��Q��� %���I�ҏm������ ���P�;�t����3� ��W���򟍟���:� ՟^�p���W����� ܯw� ���$���!�Z� ��~����=�ƿؿs� ���� ��D�߿h�� ��'ω���]��ρ�
� ��.�@�����'߈�s� ��G���k��ߏ���*� ��N���r����C� U���������8��� \���Y���-���Q��� u���������XC |�;�_�� ��B�fx %_���/� ,/�)/b/��/!/�/ E/�/�/{/�/�/(?? L?�/p??�?/?�?�? e?�?�?O�?6OHO�? �?/O�O{O�OOO�OsO �O�O�O2_�OV_�Oz_ _�_�_K_]_�_�_�_ o�_@o�_do�_ao�o 5o�oYo�o}o�o��o�o`K��y�$�REFPOS8 �1*����q� @ x +=w���=� �a��^���2���V� ߏz�������]� H������@�ɟd�Ɵ ����#���G��k�}� �*�d�ů��鯄�� ��1�̯.�g����&� ��J�ӿ忀���̿-� �Q��u�ϙ�4ϖ� ��j��ώ�߲�;�M� ����4ߕ߀߹�T��� x�����7���[��� ����P�b���� ��!���E���i��f� ��:���^����� ����eP�$� H�l��+� O�s� 2l� ���/�9/�6/ o/
/�/./�/R/�/�/ �/�/�/5? ?Y?�/}? ?�?<?�?�?r?�?�? O�?COUO�?O<O�O �O�O\O�O�O	_�O_ ?_�Oc_�O�_"_�_�_ X_j_�_o�_)o�_Mo �_qoono�oBo�ofo �o�o%�o�om X�,�P�t� ��3��W��{��� (�:�t�Տ������� ��A�܏>�w����6� ��Z��������ܟ=� (�a����� ���D��� ߯z����'�¯K�]� ��
�D�����ɿd�� ��Ϭ��G��k�� ��*ϳ���`�rϬ�� ��1���U���y��v� ��J���n��ߒ��-� �����u�`��4�� X���|������;��� _������0�B�|��� ����%��I��F �>�b�� ���E0i� (�L���/� //�S/e/ //L/�/ �/�/l/�/�/?�/? O?�/s??�?2?�?�? h?z?�?O O9O�?]O �?�OO~O�ORO�OvO �O�O#_5_�O�O_}_�h_�_�Y�$REF�POSMASK �1+����Q� �R@��_�W�WXNO  ��_�_�^MOTE�  l�TEa_CFOG ,LmgQ>T��b�QPL_RAN�GHaBQe��fOW_ER -e�`��fSM_DRYP�RG %i�%�I_�o�eTART �.�nzUME_�PRO�o�oc�T_�EXEC_ENB�  �e�iGSP�D<p~p�x�xT3DB��zRM��x�INGVERSI_ON jR��YI_AIRPUR�` DzdY��[�MIeb/LnBR� ��` ;)y�MOVH`�����EP<Ō�mz�~q �2m  >T\fT!� >W��@�R�d�v�|� X�b \�QC3�����r@�
�rA�9:�`˟�@���]������t�@�����$���@���!� d�_��_/�� $�e� ���D�������,�s�T_�PT�`Jk��eOBOT_ISOLCl�Ԡա�e��U�NAME
����A�_CATEGh�cc`�������ORD_NUM �?�hR�H705  >T������PPC_T�IMEOUT�o �x�PS232eb1�3e�s L�TEACH PENDAN/�aW����؍H_FPMa�intenanc?e Cons��|��>U"��BTNo Use؏�Ϗ�����p�#�5�D�NPOp\1a�cD�oCH_L?p4	��С	�с�!U�D1:�߃�R�PVGAIḺ1×��e�D�PACE1 {25k�� �jW܏��d�b��ի���< �U�?����������� ,�M�\�T�f�x��<� ����������1 Fgb�t�������\ �����@�Q8 f�����j� /��>/_/6/t/ �/������/� /(?I?�/�/?f?�? �?�/�/�/�/�?
?? 6O@?OlO�OdOvO�O �?�?�?�?O�O*OLO V_w_6_�O�_�_�_�_ �O�O__&_8_J_l_ voDo�o�o�o�o�o�_ o"o4o�oXozo� �d����� 0BT�x��� �ȏ�����.�,� >�P�b��������ӟ ���	���?�:�L� ^�p���4���ȟү� ���)��>�_�Z�l� ~���B�����a��� �7��L�m�h�z��� ����b�Կ�� �!��� j�W�>�lߍ߈ϚϬ� ��p���������D� e�<�N�w�ߨߺ��� �ߐ��$�.�O���� ��l������������� ���"�D�Nr� �|�������� �0R\}<�� �����, �Pr|/��/�/�/ �/�////(/:/�/ ^/�/�?�?j?�?�?�? �?O?$?6?H?Z?O ~?�?�O�?zO�O_�O _7_2ODOVOhO_�O �O�_9_�_�_o�_$o Eo@_R_d_v_�_:o�_ �_�o�o�oBo/D e`oro�o�oH�o�o ��o��=��&�O� n����h��� �'��p�]�D�r��� ������ď֏���� &���J�k�}�T�f��� ����ҟ䟖��*�4� U��j���r������� ί�����(�J�T� ��xϙϫϒϔ�޿ܿ � ����6�X�b߃� Bߘ߹ߠ��������� � �2���V�x߂����R��������� ��$RSPACE�2 25����0� ��0�B���f� �����������<�3-�?�Q�c�u� '�����F�9pNoMCE4b t���\� / {�M/n/E/�/�/�CE5����� �//5/L?�/,?�?�?pz?�?�?�/CE6�/ �/�/??�?8?j?�O �?aO�O�O�O�O_�?CE7OO%O7OIO �OmO�O�__�_�_op�_"oCo!_CE86_ H_Z_l_~_0o�_�_�o Oo�o!BWxVo�CEG 9nk� �jt
�p �  ne��� "�4�F�X�pc�hw��o p��t֏��d�� ��#�5�G�Y�k�}� s�������şכ��� ���9�K�]�o����� ������������ ���Y�k�}������������ͯ߯�� `S @LŴ� Z�6�>���µ#ϩ� �����ʜ����"�@� ��(�j�|�F�P�bߔ� �ߘߪ߼���0�B�`� �H���f�p������Ƽ
z�K�s�Y�_MODE  �nka�S :ni�# :����ovψ����
	:b�T�MP mf�`� oo�o���o�o� ��0Ef�|�CWORK_AD�q���*��!R  ��{`�?��_INTVAL�q������OPT7ION� ��!�V_DATA_G�RP 2≮��D2�P'G/#k/ V)$��/�/�/�/�/�/ ?�/??(?^?L?�? p?�?�?�?�?�? O�? $OOHO6OlOZO|O~O �O�O�O�O�O_�O2_  _B_h_V_�_z_�_�_ �_�_�_�_�_.ooRo @ovodo�o�o�o�o�o �o�o<*LN `����������8�&�\�t��$�SAF_DO_PULSq�u�l���v�CAN_TIM�p�B����R �=#h�#��~�J]]
��a!]�~ց3� `/� � 2�D�V�h����������ԟ�t#l"�2�ց�d�*�\"ԃ�O��s�t���Z>���P����B�_ @T�  �T��������T D��B�T�f� x���������ҿ��� ��,�>�P�b�_��.P�r�r�����  �;�#oV��~p���
�u��Di��S  � � �~ޅ΁��^�p� �ߔߦ߸������� � �$�6�H�Z�l�~�� ������������ � 2�D�V�h�z����������������
V� m�J\n���� ��)��*< N`r������0k�4�+�ۈ���� �////A/S/e/w/ �/�/�/�/�/�/�/? ?+?=?O?a?s?�?�? �?�?�?�?�?OO'O 9OKO]OoO�O�O�O�O �O4�O�O_#_5_G_ Y_k_}_�_��_�_�_ �_�_oo1oCo�4ћ�DЀo`jao`o`�����o�o�o �o�o�g�o�o"4 FXj|���� �����0�B�T� f�x���������ҏ䏀����,�>�P�%�� y�)�[�������Ο�� ���(�:�L�^�p� ��������ƪ��ϯ\������������	12345�678K�h!B�Q!��'Z
�����l�~��� ����ƿؿ������ %�7�I�[�m�ϑϣ� �����������!�3� E�V��yߋߝ߯��� ������	��-�?�Q� c�u���X�j����� ����)�;�M�_�q� ���������������� %7I[m� ������! 3Ei{��� ����////A/ S/e/w/�/�/Z�/�/ �/�/??+?=?O?a? s?�?�?�?�?�?�?�? �/O'O9OKO]OoO�O �O�O�O�O�O�O�O_ #_5_G_Ok_}_�_�_ �_�_�_�_�_oo1o�CoUogoyo�o�o<� i��o�o�eb_�o	�o�Cz  A��a�   �s�2��}Q��j� <�
sw_�  	�<�2�o �����|psa��l��*�<�N�`�r��� ������̏ޏ�����&�8�J�\�n����(up��(������ϟ� ���)�;�M�_�q� ��������˯ݯ��D�<��a�qYr<7�� -��q  �G�a�Ksy�D�|�q�qt  Np`����tp���� `3r D�п�A}y��6�3r��$SCR_GR�P 1?#�`�#��� 	$ ��`r Tu	 D��L�]�V��o͑�i�p�υϾ�*}�cp~��D1� D�~�c�׻��
CR�X-10iA/L� 2345678+90�p2� @уp�2�L O�3q
V14.00 l�h��R�z�s{ �ցL���;���;�� )�bq[ɏ���	�������� �2�B��G�H�L���P����G5_�B�m��D%�C6&��C3���5���B�sh�C3�����r@�
�rA�94�`�߶@��TB�  �=8B�ov�D%�C6 �L��3q�����#�T0w�i/xh7p,��?B�  B�n�l���h�ANp��  @�6p��h�@���� ?���h�Hr������h�F@ F�` �;&_Jo �����`�����`�)B�7 �}h����� ��/
/C/./g/y/@��çϙ'�/q�
�/�/��@-;��6p0?:r��F71=�V7Uv�b��?51��&@�5���3��0��23q �2�3�1�?OM�1(H4OFOO��|O��O�?�/�O�O�O�� 0�f4�3!W�O>_����ECLVL  �3q���ҷ0j7�\QL_DEFAU�L��fRW����6pxSHOT�STR�]�1�RMI�POWERFcP�2u�U[R�PWFDO��V �ZRVEN�T 1@kQkQ�S� L!DUM_�EIPJ_���j!AF_INE��!FToxnD?o�o!;´o�L��o��o!RPC_M'AIN�o�H��o4N�cVIS�I�#~�!OPCU41̜��o�!�TP�pPU�2id���!
PMON?_PROXY�5fAe�d��r2�.mfS����!RDM_S�RV��2ig����!#Rh4�3hh�H�K!
�`M{�/li7����!RLSYN�C����8����!�ROSo��4�ϟ,�!
CE�pMOTCOM-�5fk��x�!	A�CONSdy�4glg�į!A��WASRCˏ5fm쳯�!A�USB��3hn��\�!S#TM�Pv�1joK�����o̿����L_�QICE_KL ?%k� (%SVC�PRG1��=�'�2�=�B�,�3e�j�,�4��ϒ�,�5�Ϻ�,�6����,�7�
�,�]�$M�H�9U�Z�)�� ��,�/Ϫ�,�W���,� ���,���"�,���J� ,���r�,�ߚ�,�G� ��,�o���T����T� ��:�T���b�T��� T�8��T�`���T��� T���*T���RT�  �z|�(����,�� %��
��2V Aze����� ��//@/+/d/O/ v/�/�/�/�/�/�/? �/*?<?'?`?K?�?o? �?�?�?�?�?O�?&O OJO5OnOYO�O�O�O �O�O�O�O_�O4__�F_j_U_�_ �_DE�V i��UT1:����4�TGRP 2D�e�P!�bx 	�� 
 ,�P �Q�_o�T.o@o'odo Ko�o�o�o�o�o�o�o �o�o<#`rY �}{�U���yo� �$��H�/�l�~�e� ����Ə؏����� � 2��V��z���C�� ��C�ܟß ����6� �Z�A�S���w����� د�ѯ�e���D��� h�O�������¿��� ��߿��@�R�9�v� ]Ϛρϓ���'���� ��*��N�5�G߄�k� �ߏ����������&� 8��\�C����϶� m����������4�F� -�j�Q���u������� ����B��7 x/������ �,P7t� m�����/[ (/:/!/^/E/�/i/{/ �/�/�/�/ ??�/6? ?Z?l?S?�?w?�?�? /�?�?O OODO+O hOzOaO�O�O�O�O�O �O�O__@_R_9_v_��Yd �Xzh9�6T 	 �A��:��A36|=>����h�@�- ��Z�P�G�A=���?�&%�H��@�������]B���A�|�����?����§=������]@��}����AÖ�@��h�����AZ��Y%P�ROVA�_Xo���la�Qle|o�g�to�o�o�o�o�o y%�Yo'  �o�o J�n���
� .�"��2�4�F�|� j����Ǐ������ ��.�0�B�x����� ޏh�ҟ������� *�����w���P����� ί�����X�=�|� �p��������ʿ�� �0��T�޿H�6�l� Z�|Ϣϐ������,� �� ��D�2�h�V�x� ������ߎ������ 
�@�.�d�ߋ��T� v�P��������<� ~�c���,��������� ������V�;z� n\������ .R�F4jX �|���*� //B/0/f/T/�/� �/�z/�/v/�/?? >?,?b?�/�?�/R?�? �?�?�?�?OO:O|? aO�?*O�O�O�O�O�O �O�O_TO9_xO_l_ Z_�_~_�_�_�__�_ o�_�_�_2ohoVo�o zo�o�_�oo�o
�o .dR��o� �ox������ *�`�����P����� ޏ̏����h���_� ��8���������ڟȟ ��@�%�d��X��h� ��|�����֯���<� Ư0��T�B�d���x� ���տ������,� �P�>�`φ�ȿ��� v��������(��L� ��s߅�<�^�8ߦ��� �� ���$�f�K��� ~�l���������� >�#�b���V�D�z�h� �����������:��� .R@vd��� ���* N<r���b� ^�/�&//J/� q/�:/�/�/�/�/�/ �/�/"?d/I?�/?|? j?�?�?�?�?�?�?<? !O`?�?TOBOxOfO�O �O�OO�O�O�O�O�O _P_>_t_b_�_�O�_ �O�_�_�_oooLo :opo�_�o�_`o�o�o �o�o�o H�oo �o8������ �PvG�� �z�h� �������(��L� ֏@�ҏP�v�d����� �� ��$�����<� *�L�r�`���؟���� ���ޯ��8�&�H� n�����ԯ^�ȿ��� ڿ���4�v�[�m�$� F� ώ��ϲ������ N�3�r���f�T�v�x� ���߮���&��J��� >�,�b�P�r�t��� ����"����:�(� ^�L�n��������� ���� 6$Z�� ���J�F��� �2tY�"� z�����
/L 1/p�d/R/�/v/�/ �/�/�/$/	?H/�/<? *?`?N?�?r?�?�/�? �?�?�?�?O8O&O\O JO�O�?�O�?pO�O�O �O�O�O4_"_X_�O_ �OH_�_�_�_�_�_�_ �_0or_Wo�_ o�oxo �o�o�o�o�o8o^o/ nobP�t�� ��4�(��8� ^�L���p����͏� �� ��$��4�Z�H� ~������n�؟Ɵ�� � ��0�V���}��� F�����ԯ¯���� ^�C�U��.��v��� ��п����6��Z�� N�<�^�`�rϨϖ��� ���2ϼ�&��J�8� Z�\�nߤ�����
ߔ� ����"��F�4�V�� �ߣ���|��������� ��B���i���2��� .�����������\� A��
tb��� ���4X�L :p^���� �0�$//H/6/l/ Z/�/��/�/�/�/|/ �/ ??D?2?h?�/�? �/X?�?�?�?�?�?O 
O@O�?gO�?0O�O�O �O�O�O�O�O_ZO?_ ~O_r_`_�_�_�_�_ �_ _F_oV_�_Jo8o no\o�o�o�o�_�oo �o�o F4jX ��o��o~��� ��B�0�f����� V������ҏ���� >���e���.������� ����Ο�F�+�=��� ��^���������ܯ ��B�̯6�$�F�H� Z���~�����ۿ��� ���2� �B�D�Vό� ο���|�����
��� .��>ߔϺϋ���d� �߬��������*�l� Q�������� �����D�)�h���\� J���n���������� @���4"XF| j������ �0TBx�� �h�d�/�,/ /P/�w/�@/�/�/ �/�/�/?�/(?j/O? �/?�?p?�?�?�?�? �? OB?'Of?�?ZOHO ~OlO�O�O�OO.O�O >O�O2_ _V_D_z_h_ �_�O�__�_�_�_o .ooRo@ovo�_�o�_ fo�o�o�o�o* N�ou�o>��� ��� �&�hM��u��p�$SERV�_MAIL  ʌu����ql�OU�TPUTw���p@l�RV �2E�i��  �(�R�ޏl�SAV�E����TOP10� 2F�� d o6�� (� F�X�j�|�������ğ ֟�����0�B�T� f�x���������ү� ����,�>�P�b�t� ��������ο���0�(�:��YP�����FZN_CFG ;G����t����r�GRP 2�H|�	� ,B �  A���qD;�� B���  B�4�sRB21��HELLu�I��ˀ̏��%�4�%RSR4�5�G� ��kߤߏ��߳����� ��"��F�1�j�U�������  �h�%����������	���p������w��2�pd�	�����HK 1J�� "����������� ����61CU~ y��������?OMM K��5���FTOV_EN�Bw�h��HOW_?REG_UIU���IMIOFWDL� L$�ŊWAITR��²��v����TIMv���VAv���_UNITQ &��LCoTRYv��l�MB_HD�DN 2M�� ����u� ��/� �/�/�/�/�/"??+?(X?^2r!Eu�N�ɧ��Y�p3��O|; �����<�u>Ak����X�px��,��?�  �?d�;Ʉi�u�i�彌p6�9�q<, � :�  =@=7���JËtG@�`G�MO�N_ALIAS k?e$ǀhe=� �O�O�O�O�J�O__ /_A_�Oe_w_�_�_�_ X_�_�_�_oo�_=o Ooaoso�o0o�o�o�o �o�o�o'9K�o o����b�� ��#��G�Y�k�}� ��:���ŏ׏鏔�� �1�C�U� �y����� ����l����	��-� ؟Q�c�u���2����� ϯ�󯞯�)�;�M� _�
���������˿v� ���%�7��[�m� ϑ�<ϵ��������� ��!�3�E�W�i�ߍ� �߱����߀����� /���@�e�w���F� �����������+�=� O�a�s���������� ����'9��] o���P��� ��5GYk} (������/ /1/C/�g/y/�/�/ �/Z/�/�/�/	??�/ ??Q?c?u?�?2?�?�? �?�?�?OO)O;OMO��?qO�O�O�O�ObC��$SMON_DE�FPROG &�����A� &*SYS�TEM*�O�O�BR�ECALL ?}~�I ( �}kO@O_a_s_�_�_�_ =_ �_�_�_oo(o�_Lo ^opo�o�o�o9o�o�o �o $�oHZl ~��5���� � ��D�V�h�z��� ��1�ԏ���
�� ��@�R�d�v�����-� ��П�����*��� N�`�r�������;�̯ ޯ���&���J�\� n�������7�ȿڿ� ���"ϵ�F�X�j�|� �Ϡ�3���������� ߱�B�T�f�xߊߜ� /������������ +�P�b�t����=� ��������(���L� ^�p�������9����� �� $��HZl ~��5����  �DVhz� �1����
// �@/R/d/v/�/�/-/ �/�/�/�/??*?�/ N?`?r?�?�?�?;?�? �?�?OO&O�?JO\O nO�O�O�O7O�O�O�O �O_"_�OF_X_j_|_ �_�_3_�_�_�_�_o o�_BoTofoxo�o�o /o�o�o�o�o�o +Pbt���= �����(��L� ^�p�������9�ʏ܏�� ��$����$S�NPX_ASG �2P���J��� P 0� '%R[?1]@1.1+���?���%u���M��� ȟ{������"���� X�;�M�����u�����abX��诛�ݯ �q�B���7�x�+�m� ����ҿ�ǿ���� >���b�E�WϘ�[����ϸ�&��Ϫ���-� ��Q��F߇�:�|߽� ������������M� ��q�T�f��jߜ������4������� >���b��W���K��� ��������( ^���ew�{�� ���H�= ~1�U���� /A2/D/'/h/�]/ �/�/�/��/�/�/�/ .??R?5?G?�?k?}?��?�/�?�?�?O�� OGOJ/<O}O�?�O�? �O�O�O�O_�O1__ &_g_J_\_�_�_�_�_�_�_�X%�_'oZOo ]o@o�o�_o�o�O�o��o�o�oGʨn�7x+m����~���ko�>�!��=�PARAM �QJ�T� ��	��P�e�������� ��=�O�FT_KB_CF�G  �tQ�:�O�PIN_SIM  J���������[�RVNORDY_DO  ���ǅ/�QSTP_DSBێ��s�Wx�[�SR Rމ� � &��OS2�  ORT�Wy��u��TM_CTL� 3Sޅ��  p%|�	��-� ��B�Q�[t��|���1� C�^sށ_������ ��˯�^�p��%�7� I�ʿܿ�����6��H�Z���χ��GR�Pۈ�p���OP_?ON_ERR<��ƿPTN ��D��RING_�PRM��N�VCNT_GP 2Tޅ:����x 	��`��_pN߇�r߫ߊ�VDL5Т�1Uj����� ��������
��.�U� R�d�v������� ������*�<�N�`� r��������������� &8J\n� ������� "4Fmj|�� �����/3/0/ B/T/f/x/�/�/�/�/ �/�/�/??,?>?P? b?t?�?�?�?�?�?�? �?OO(O:OLO^O�O �O�O�O�O�O�O�O _ _$_K_H_Z_l_~_�_ �_�_�_�_�_oo o 2oDoVohozo�o�o�o �o�o�o�o
.@ Rdv����� ����*�<�c�`��r�����������PR�G_COUN��r͔����ENB���M���_UP�D 1V��T  
Ϗ&�b�t����� ����Ο�����?� :�L�^���������ϯ ʯܯ���$�6�_� Z�l�~�������ƿ� ����7�2�D�V�� zόϞ���������� 
��.�W�R�d�vߟ� �߬߾��������/� *�<�N�w�r���� ���������&�O� J�\�n����������� ������'"4Fo j|��������،_INFO� 1WP��6�X	 ;����?>�?���>P`=f�_3;3����/ܛ^n�jQ��]=.^������zC3ҍ�����@�, A�����`�9@��z�=�@ �>/ȝ ����CD25D�4�1Ca������<&/�8'�YSDEBU)G��Q��%d�a SP_PASS���B?s+LOG �XMZ�  z%�!?���%�,  �5�%UD1:\�$3�"o_MPC�/ �$(�",?�,�(2�/2?SAV Y�)��؉�!(:�(SV�`;TEM_TIM�E 1Z�'[�� 0  V��K�2?�3�3MEM�BK  P�5��� �/5OGOWLX�|6�� @WO$��yO�O�LrO�O,�Jn! �@�1_ (_:_L_�3d_v_�_�_�_�_�_ ��_�_o o,o>oPoboto�o��e�o�o�o�o�o &8J\n�����������5S!K@H�� K �_��q�eGM�`T�L�  D�O�� �-�H�O���O�H	A�_��E�W�%`Q_��  ���H�M�lȟڟ ߏ ����B��7�I�[�m��%U�����o˯!{ӯ��	��-�?� Q�c�u���������Ͽ�����)�9T1SVGUNSP����# 's%�D�2�MODE_LIMG [�9w"@�2M��m�\�-?�ABU�I_DCS _3�s!#@�������C 2������C *���=� 
C�,=�@��W�(�7X��,��EDIT `����&9�  E�;���CZ  C�$H��SCRN �a�-���0��-,)� �cD��	0OG b���؅6����SK_OPTI�ONh Iw!��_D�I� ENB  ��s%��BC2_G_RP 2d���� X�ϺD�PC8����a?%�����CFI��f��&=��(?C� o�������������� �� 9$IoZ �~������ �5 YD}h� �������/+/ =/�a/L/q/�/�/�/ ��3��/@� �/?�/ (??L?:?p?^?�?�? �?�?�?�?�?O O6O $OFOlOZO�O~O�O�O �O�O�O�O�O2_X�� F_X_v_�_�__�_�_ �_�_�_o*o<o
o`o No�oro�o�o�o�o�o �o&J8n\ ~������� � �"�4�j�X���D_ ����֏���x��� .�T�B�x�����j��� ���ҟ�����,� b�P���t�����ί�� ޯ��(��L�:�p� ^�������ʿ��� ��6�H�Z�ؿ~�l� �ϴϢ��������� � �D�2�h�V�x�zߌ� �߰�����
���.�� >�d�R��v����� ��������*��N�� f�x�������8����� ��8J\*� n������� "F4jX�| �����/�0/ /@/B/T/�/x/�/d� �/�/�/??�/>?,? N?t?b?�?�?�?�?�? �?O�?(OO8O:OLO �OpO�O�O�O�O�O�O �O$__H_6_l_Z_�_ ~_�_�_�_�_�_o�/ &o8oVohozo�_�o�o �o�o�o�o
�o@ .dR�v��� ����*��N�<� ^���r�����̏���� ޏ ���J�8�n�$o ������ȟڟX������4�"�X�B�v��$�TBCSG_GR�P 2gB���  �v� 
 ?�  �� ����ׯ�������1���U�g�z���i��_d�H��?v�	 HA���e��>���>f���\e�AT��A ���пܸ�����G��?L��Ʋpܿ޾�;ff�������v�򾺠$�l�@��R����ff>�33��e�~�B˿m��J�����Ɍ�϶�҃�H��B����B��϶�K�E�K�j�}� H�Zߨ��ߐߢ�������ؐ6�	V3�.00��	cr;xl�	*X�P�u���[���H���� q��p��  O��Cp�����z�J2ʁ�k�����#�	 @����8�J�\�n��������������CFoG mB���Y ��#����9#�/�/U (���s���� ��*N9r ]������� /�8/#/\/G/�/�/ }/�/�/�/�/�/?3 ��?.?@?�/s?^?�? �?�?�?�?�?�?O'O 9OKOOoOZO�O~O�O �Ov�b��O>��O __ H_6_l_Z_�_~_�_�_ �_�_�_o�_2o oVo Dofohozo�o�o�o�o �o�o
,R@v d�������� ��<�*�`�N���r� ����̏ޏ������ 8�&�\�n�����L��� ��ڟȟ����4�"� X�F�|�j�������֯ į�����B�0�R� T�f����������ҿ ����>��V�h�z� $ϪϘϺϼ������ (��L�^�p߂�@ߦ� ���߸��� ��$��� 4�Z�H�~�l����� �������� ��D�2� h�V���z��������� ��
��.>@R �v������� ��N<r`� �����//� $/J/8/n/\/�/�/�/ �/�/�/�/?�/ ?F? 4?j?X?�?|?�?�?�? �?�?O�?0OOTOBO xOfO�O�O�O�O�O�O �O__*_,_>_t_� �_�_�_Z_�_�_�_o o:o(o^oLo�o�o�o �ovo�o�o �o6 HZ&�~�� �����2� �V� D�z�h��������� ����
�@�.�d�R� t����������П� ��_0�B��_����r� ����̯��ܯ��&� 8�J�����n����� ȿڿ�����"��2� 4�F�|�jϠώ��ϲ� ��������B�0�f� Tߊ�xߚߜ߮����� ���,��P�>�`�� t��$�V������� ��L�:�p�^����� ���������� " $6l~��\� ���� 2 hV�z���� �
/�.//R/@/v/ d/�/�/�/�/�/�/�/ ??<?N?��f?x?�? 4?�?�?�?�?�?�?O 8O&O\OnO�O�OPO�O�O�O�O�O�N  $P(S (V<_(R��$TBJOP_�GRP 2n�E��  �?���C(R	�TR[Spb\��@��X  �(U�P �, � ��P^(S @$P?�Q	 �A����U?C�  DBW�Q��Q>tP>\?�`�UaG�:��o�];ߴAgT���U�QA�:c��UKoVg�_�_>�Q��\)?���f8�Q��Q�RL��>y�.`$P;iG,b��gAp:`�`Do�oA�ff�eto�T�`xr'~:VM�,b���`Qt<om(U@�;�R�uCр�Q��Q�u�t�b�e�ff��u:�6/�q?�{33�uB   �q �����r�a�d�}^<�:�S��~��px}�����@��H���$��x-q�p�u=�`<�#�
(v�QtP;/��ڨ�?��P�B�
��%�0i�U0�fw X�B�P�~�����D�Ο �ҟ���?��ԟ^��x�b�p���ϯ(SC��(V���U	V3�.00yScrxl�T*��T#Q��at3� F�� H�H F6�� F^ F��� F�f F�� G� G5� G<
 G^]� G� G����G�*�G�S� G�; G���C�Dup��E[�� E� F(� F-� FU`� F}  F�N� F� F��� Fͺ F�� F�V G�� Gz Ga� 9ѷ챸�HD �d�2_�*�(V�.� ��U��F^ED_TCH qb[�)�0�
(  ��u$Pd$%�����(TB�����C��U���STPARS  �X��TPHR �A�BLE 1rbYC L����C� �0#�������'W/Q*��	��
����Zժ(Q������N7�RDIB�lQY�@k�}ߏߡ߳��O#�5�?�Q�c�u��;�S!�jS ��H�Z�l�~� ��������������  2DVhz�� G] �$�kRX��	���� ����߼���������;��NUM  V�ElQ�P0P� W��;�_CFGG s�[�Q@TP�IMEBF_TT�&�V����VER��Q&�R 1=tJ� 8��(R�#Pc! �@�   K/]/o/�/�/�/�/�/ �/�/�/?#?5?G?Y? k?}?�?�?�?�?O�?��?OO1OCN� WOiOCN!S�O�O�O�O �O�O�O_"_4_F_X_ j_|_�_�_�_�_�_�_ �_oo0oBoTofj0$�_�&@'%��L�IF u���"!��d"!�d(�D�
����@pd� d	}��`SC�RN v� �IOx_CUR ew����	)D��O{PREV �xc}�VtS��2y�c{ xDO��) ��}g1���m�b�l�d��qMI_CH�AN� '% e�D_BGLVL����e�ETHERADW ?*����.��0Ā:eǀ4:�7d:bc:db� ďc׏dd�d�e��ROUT !��!�8�w�h�?SNMASK��'#~��255.v���t��������OOLOFS_DI&��՚�ORQCTRL zJۓ�/��T�:�L�^�p��� ������ʯܯ� �� $�6�H�Z�j����|����}�PE_DET�AI��ۚPGL_�CONFIG ������/c�ell/$CID?$/grp1��+� =�O�a�sώ���� ���������χ��.� @�R�d�v�ߚ߬߾� �����߃ߕ�*�<�N� `�r��������� �����&�8�J�\�n� ���!������������}��FXj|@��s������� �!3EW��{ �����d�/ ///A/S/e/��/�/ �/�/�/�/r/??+? =?O?a?�/�?�?�?�? �?�?�?�?O'O9OKO ]OoO�?�O�O�O�O�O �O|O_#_5_G_Y_k_ }__�_�_�_�_�_�_ �_o1oCoUogoyoo �o�o�o�o�o�o	���User �View �}}�1234567890:L^p����t ��� y2 -y�o��"�4�F�X���'r3�����ʏ@܏� �_�!��~4�� Z�l�~��������՟�~5I�� �2�D�V�h�ǟ���~6��¯ԯ����
��{�=��~7 ��v���������п/���~8e�*�<�N�`��rτ�㿥ϫ� �lCamera+z!������ �2�D�"E��n߀ߒ�8��߾����������  ���y��V�h�z�� ���W�������C��@.�@�R�d�v������ �����������
 ��@Rd����� �������H�y. @Rdv�/�� ��//*/</N/ ���"���/�/�/�/ �/�/�?,?>?�/b? t?�?�?�?�?c/�Ű� Q?OO*O<ONO`O? �O�O�O�?�O�O�O_ _&_�?��d��Or_�_ �_�_�_�_sO�_oo __8oJo\ono�o�o9_ ���)o�o�o& 8�_\n��o��@�����o�g9� ?�Q�c�u�����@�� ϏᏈ��)�;�M�(_�q� �	��0���� ��П������*�<� N���r���������̯ s�������p�%�7�I� [�m��&�����ǿ� ����!�3�E���� 9�ܿ�ϣϵ������� ���!�3�~�W�i�{� �ߟ߱�Xϒ���H��� �!�3�E�W���{�� �������������� ������i�{����� ����j�����V�/ ASew�0���}+  ���/�� Sew����� ������;�A/S/ e/w/�/�/B�/�/�/ ./??+?=?O?a?-  )�?�?�? �?�?�?�?O O2ODOVK   f?}Oh? VOx:�O�O�O�O__ )_;_M___q_�_�_�_ �_�_�_�_oo%o7o Io[omoo�o�o�o�o �o�o�o!3EW i{������A}
 (  �0( 	 ��� 2� �V�D�z�h��������ԏ�����J�J ̰/a�s��� �/����͟ߟ��
# P�-�?�Q���u����� ����ϯ����^� ;�M�_�q�����ܯ�� ˿ݿ$���%�7�I� [Ϣ����ϣϵ����� �����!�3�z�W�i� {��ϟ߱��������� @��/�A��e�w�� ���������� `�=�O�a�s������� ������&�'9 K]�������� ���#j|Y k}������ �B/1/C/�g/y/ �/�/�/�//�/�/	? P/-???Q?c?u?�?�/ �/�?�?�?(?OO)O ;OMO_O�?�O�O�O�? �O�O�O__%_lOI_ [_m_�O�_�_�_�_�_8�_2_�@ bo�,o>ocg�p���"frh:\tp�gl\robot�s\crxxa10�ia_l.xml �_�o�o�o�o�o�o0+=O��Pu �������� �)�;�RL�q����� ����ˏݏ���%� 7�N�H�m�������� ǟٟ����!�3�J� D�i�{�������ïկ �����/�F�@�e� w���������ѿ��� ��+�B�<�a�sυ� �ϩϻ��������� '�>�8�]�o߁ߓߥ� �����������#�5�:Wh�Q ob`�<< `` ?�5�x�5�p����� �������,��$�F� t�Z�|����������������(6V<P(��$TPGL_OUTPUT �@Q�@QS   h}������ �1CUgy �������	/�/hX��- cel�l/floor/�wall 8901234567P/ b/t/�/�/�%6R- �/ �/�/�/??�/�/J?@\?n?�?�?�?<7}�? �?�?�?	OO�?�?QO cOuO�O�O�OCO�O�O �O__)_�O7___q_ �_�_�_?_Q_�_�_o o%o7o�_Eomoo�o �o�oMo�o�o�o! 3�o�oi{��� �[����/�A� �O�w���������W� i�����+�=�O�� ]���������͟e�۟���'�9�K��2 $$%/�� ������ׯɯ���� �C�5�g�Y���}��� ��ӿſ�����?�@1�c�Uχ�yϫ�}S�����������0�@�Z�T�f�`� ( 	 �ϛ߉߿߭� ���������+�a� O��s�������� ���'��K�9�o�]�������������3&�  <<�� "4m [mG� �-*���� �Rd�h�4 ����//v / N/�:/�/�/p/�/�/ */�/??�/8?J?$? V?�?�/�/�?�?b?�? �?�?�?4OFO�?jO|O OhO�O�O�O�O�OXO _0_�O_f_x_R_�_ �__�_�_�_�_o,o o4obo�_Jo�o�oDo �o�o�o�oto�oL ^�oj�n��� :����H�Z�4� ~����x�Ə`����� ��2�D���,�z��� &�����Ο��V�h� .�@�ڟH�v�P�b��� ���������*����`�r�)WG?L1.XML0ߧ���$TPOFF_�LIM 	 =�����N_S]V��  7�Ϻ�P_MON ��Ѵ=�=�2���STRTCHK' �϶�ϸ��VTCOMPAT��n�ӶVWVAR� ����� KE� ��=�����_DEFPR�OG %3�%�ROS�߱�_DISPLAYİ�3���INST_M�SK  +� ~�INUSERd���LCKm�4�QU?ICKMEN���oSCRE��~o�tpscԠm�����ϲ��_��S�Tb�ϹRACE_�CFG ������	��
?�~,�HNL 2�����P�� ������������.�I�TEM 2�p�� �%$1234?567890W�i�  =<a�������  !������ k�����U�y�9K ��a�����	�- ���u���� 7����)�M _q��A/g/y/� �///%/�/�/[/? -?�/9?�/�/�?�/�? ?�?�?E?�?i?�?DO �?_O�?oO�O�OO�O /OAOSO�OwO#_I_[_ �O_�O�O_�_�_=_ �_os_o�_�_ro�_ �o�_�o�o'o�oKo]o &�oA�oQw�o�o �o+5�Y�+� =��a����c�� ��ߏ�U���y����� !�o�ӏ����	���-� ?��c�#���G�Y��� o��3����ׯ;�� ����+�����˯E� ﯛ���ӿ7���[�m� ��ϵ�uχ�뿓� �!���E��i�)�;�@��Q����Ϟ�*�S6���<���  ��� H�����
� �-��Q����UD1:\^������R_GRP 1��D�� 	 @@������������#���3�J�X���^��m�����?�  ���������� ;)KM_�� �����7�	q�K]��SC�B 2���  �������//�'/9/��UTORIAL ���E�/���V_CONFIG ���C���A���/�-OUTPUT� ���� ���/3?E?W?i?{?�? �?�?�?�?�?�?O�!  ?3OEOWOiO{O�O�O �O�O�O�O�O_O/_ A_S_e_w_�_�_�_�_ �_�_�_o_+o=oOo aoso�o�o�o�o�o�o �o&o9K]o �������� �"5�G�Y�k�}��� ����ŏ׏����� 1�C�U�g�y������� ��ӟ���	��,�?� Q�c�u���������ϯ ����(�;�M�_� q���������˿ݿ� ��$�7�I�[�m�� �ϣϵ���������� !߽/�%?_�q߃ߕ� �߹���������%� 7�*�[�m����� ���������!�3�D� W�i�{����������� ����/AR�e w������� +=Nas� ������// '/9/J]/o/�/�/�/ �/�/�/�/�/?#?5? G?X/k?}?�?�?�?�? �?�?�?OO1OCOT? gOyO�O�O�O�O�O�O �O	__-_?_POc_u_ �_�_�_�_�_�_�_o o)o;oMo^_qo�o�o �o�o�o�o�o%�7I,���� hzdqS�H��� ���#�5�G�Y�k� }�����Toŏ׏��� ��1�C�U�g�y��� ������ӟ���	�� -�?�Q�c�u������� ��ϯ����)�;� M�_�q���������˿ ݿ���%�7�I�[� m�ϑϣϵ�ƿ���� ���!�3�E�W�i�{� �ߟ߱���������� �/�A�S�e�w��� �����������+� =�O�a�s��������� ������'9K ]o������� ��#5GYk�}�����$T�X_SCREEN� 1�|u�dp�}ipn�l/�gen.htm�/'/9/K/]/�� Panel� setupa,}�/pip/rm�i_log.txta/�/�/�/�/�/q �RMI_LOG�/ }�?>?P?b?t?�?�?,?"?�?�? �?OO)O�?MO�?qO �O�O�O�O�OBOTO_ _%_7_I_[_�O _�O �_�_�_�_�_�_t_!o �_EoWoio{o�o�oo (o�o�o�o/�o �o�ow������H��UALRM_MSG ?��� ��
*�<� m�`�����������؏�ޏ��3�&�W��S�EV  ����	�ECFG ���  ��@�  A�� �  B��
  X�������"�4� F�X�j�|����������GRP 2���� 0�	 ?��1�>��q�(�P���i��?� ��^�I_BB�L_NOTE ����T��#l�������DEFPR0?%� (%K�r�� �`�����ROS2 ��x�ƿ�ֿ���3���W�B�{ύ��FK�EYDATA 1y���p ��� ������6�0�� �2��,(��c���Qߎ�u�CAN�CEL����(	P�REV STEP��n�EXT���{�INISH�F�}��ORE INFO G�J�������� �������;�M�4�q��X����� ���/frh/gui�/whiteho?me.png������
.�/Se�w���</F�RH/FCGTP�/wzcancel����!3>=�
prev�m����<�	next\�//'/9/��wzfinish�w/�/�/�/�/N-infof/�/	?? -???:c?u?�?�?�? �?L?�?�?OO)O;O MO�?qO�O�O�O�O�O ZO�O__%_7_I_�O m__�_�_�_�_�_h_ �_o!o3oEoWo�_{o �o�o�o�o�o���o /ASelo�� ����r��+� =�O�a��s������� ͏ߏ񏀏�'�9�K� ]�o���������ɟ۟ �|���#�5�G�Y�k� }������ůׯ��� ���1�C�U�g�y�� ������ӿ���	Ϙ� -�?�Q�c�uχ�ϫ� ��������ߔ��;� M�_�q߃ߕ�$߹��ߠ������� �}������I�@[�m�E���{�,�� ��������,��P� 7�t���m��������� ����(:!^E �i�����  �o6HZl~� �ߴ����/ / �D/V/h/z/�/�/-/ �/�/�/�/
??�/@? R?d?v?�?�?�?;?�? �?�?OO*O�?NO`O rO�O�O�O7O�O�O�O __&_8_�O\_n_�_ �_�_�_E_�_�_�_o "o4o�_Xojo|o�o�o �o�oSo�o�o0 B�ofx���� O����,�>�P� 't���������Ώ� ���(�:�L�^�� ��������ʟܟk� � �$�6�H�Z��~��� ����Ưد�y�� � 2�D�V�h��������� ¿Կ�u�
��.�@� R�d�v�ϚϬϾ��� ���σ��*�<�N�`� r�ߖߨߺ������� ��&�8�J�\�n�� ������������ "�4�F�X�j�|���e�����e����������������,�B�fM� ������� >P7t[�� �����/(// L/3/p/�/a��/�/�/ �/�/ ?�$?6?H?Z? l?~?�??�?�?�?�? �?O�?2ODOVOhOzO �OO�O�O�O�O�O
_ _�O@_R_d_v_�_�_ )_�_�_�_�_oo�_ <oNo`oro�o�o�o7o �o�o�o&�oJ \n���3�� ���"�4��X�j� |�������A�֏��� ��0���T�f�x��� �������/����� ,�>�E�b�t������� ��ί]����(�:� L�ۯp���������ʿ Y�� ��$�6�H�Z� �~ϐϢϴ�����g� ��� �2�D�V���z� �ߞ߰�������u�
� �.�@�R�d��߈�� �������q���*� <�N�`�r�������� �������&8J \n�������h��Ր �Ր���);M%o�[,m/�e/ ���/�0//T/ f/M/�/q/�/�/�/�/ �/???>?%?b?I? �?�??�?�?�?�?џ O(O:OLO^OpO�O �O�O�O�O�O _�O$_ 6_H_Z_l_~__�_�_ �_�_�_�_�_ o2oDo Vohozo�oo�o�o�o �o�o
�o.@Rd v������ ���<�N�`�r��� ��%���̏ޏ���� ��8�J�\�n������� 3�ȟڟ����"��� F�X�j�|�����/�į ֯�����0�OT� f�x���������ҿ� ����,�>�Ϳb�t� �ϘϪϼ�K������ �(�:���^�p߂ߔ� �߸���Y��� ��$� 6�H���l�~���� ��U������ �2�D� V���z����������� c���
.@R�� v������q *<N`�� �����m//@&/8/J/\/n/E�p+��E������/�/�-�/�/�/�&, �?"?�?F?-?j?|?c? �?�?�?�?�?�?�?O 0OOTO;OxO�OqO�O �O�O�O�O_�O,__ P_b_A��_�_�_�_�_ �_�oo(o:oLo^o po�_�o�o�o�o�o�o }o$6HZl�o ��������  �2�D�V�h�z�	��� ��ԏ������.� @�R�d�v�������� П������*�<�N� `�r��������̯ޯ �����8�J�\�n� ����!���ȿڿ��� ϟ�4�F�X�j�|ώ� ��w_���������� %�B�T�f�xߊߜ߮� =���������,�� P�b�t����9��� ������(�:���^� p���������G�����  $6��Zl~ ����U��  2D�hz�� ��Q��
//./ @/R/�v/�/�/�/�/ �/_/�/??*?<?N? �/r?�?�?�?�?�?�?ڵ��;������	OO-MOOOaO;F,M_�OE_�O�O �O�O�O_�O4_F_-_ j_Q_�_�_�_�_�_�_ �_�_ooBo)ofoxo _o�o�o�o�o���o ,>P_?t�� ����o��(� :�L�^���������� ʏ܏k� ��$�6�H� Z�l���������Ɵ؟ �y�� �2�D�V�h� ��������¯ԯ��� ���.�@�R�d�v�� ������п������ *�<�N�`�rτ�Ϩ� ��������ߑ�&�8� J�\�n߀�ߤ߶��� ��������o4�F�X� j�|��߲������� ������B�T�f�x� ����+��������� ��>Pbt�� �9���( �L^p���5 ��� //$/6/� Z/l/~/�/�/�/C/�/ �/�/? ?2?�/V?h? z?�?�?�?�?Q?�?�? 
OO.O@O�?dOvO�O �O�O�OMO�O�O__�*_<_N_%�P[�>%����y_�_ �]u_�_�_�V,�oo �o&ooJo\oCo�ogo �o�o�o�o�o�o�o 4XjQ�u� ������0�B� !�f�x����������O �����,�>�P�ߏ t���������Ο]�� ��(�:�L�۟p��� ������ʯܯk� �� $�6�H�Z��~����� ��ƿؿg���� �2� D�V�h����Ϟϰ��� ����u�
��.�@�R� d��ψߚ߬߾����� �߃��*�<�N�`�r� ����������� �&�8�J�\�n���W� �������������" 4FXj|�� �����0B Tfx���� ��//�>/P/b/ t/�/�/'/�/�/�/�/ ??�/:?L?^?p?�? �?�?5?�?�?�? OO $O�?HOZOlO~O�O�O 1O�O�O�O�O_ _2_ �OV_h_z_�_�_�_?_ �_�_�_
oo.o�_Ro�dovo�o�o�o�o����k�������o�o}�o/Av,-�r%��}�� ����&��J�1� n���g�����ȏڏ�� ���"�	�F�X�?�|� c�������֟���� �0�?oT�f�x����� ����O������,� >�ͯb�t��������� K�����(�:�L� ۿpςϔϦϸ���Y� �� ��$�6�H���l� ~ߐߢߴ�����g��� � �2�D�V���z�� �������c���
�� .�@�R�d�������� ������q�*< N`������� ��ǟ&8J\ nu������ ��"/4/F/X/j/|/ /�/�/�/�/�/�/�/ ?0?B?T?f?x?�?? �?�?�?�?�?O�?,O >OPObOtO�OO�O�O �O�O�O__�O:_L_ ^_p_�_�_#_�_�_�_ �_ oo�_6oHoZolo ~o�o�o1o�o�o�o�o  �oDVhz� �-����
���.�0�����Y�k�}�U�������,��⏕�� �*�<�#�`�G����� }�����ޟ�ן��� 8�J�1�n�U���y��� ȯ���ӯ�"�F� X�j�|������Ŀֿ �����0Ͽ�T�f� xϊϜϮ�=������� ��,߻�P�b�t߆� �ߪ߼�K������� (�:���^�p���� ��G����� ��$�6� H���l�~��������� U����� 2D�� hz�����c �
.@R�v �����_�/ /*/</N/`/7��/�/ �/�/�/�/�??&? 8?J?\?n?�/�?�?�? �?�?�?{?O"O4OFO XOjO�?�O�O�O�O�O �O�O�O_0_B_T_f_ x__�_�_�_�_�_�_ �_o,o>oPoboto�o o�o�o�o�o�o�o (:L^p�� ���� ���6� H�Z�l�~������Ə ؏������2�D�V��h�z������$UI�_INUSER � �������  �����_MENHI�ST 1���  (ΐ�w '/SOFT�PART/GEN�LINK?cur�rent=men�upage,71,1 15ޟS�e�$w��)�*�1��=��ůׯ�������37=��Z�l�~����1�163¯ۿ�����+�*��2�8<�30�c�uχ��(�:�3˿�����ߧϹ�7�4��f�xߊߜ�#�=�G�22������$���*��7�B�T� f�x���� >��� ����	��-���Q�c� u�������:������� );��_q� ���H�� %7�[m�� ��V��/!/3/ E/0�i/{/�/�/�/�/ �/��/??/?A?S? �/w?�?�?�?�?�?`? �?OO+O=OOOaO�? �O�O�O�O�O�OnO_ _'_9_K_]_�O�_�_ �_�_�_�_�_|_o#o 5oGoYokoV/to�o�o �o�o�o�o�_1C Ugy���� ����-�?�Q�c� u��������Ϗ�� ���)�;�M�_�q��� �����˟ݟ��� ��7�I�[�m����|o *�ǯٯ����!�$� E�W�i�{�����.�ÿ տ�����/Ͼ�S� e�wωϛϭ�<����� ����+ߺ�O�a�s� �ߗߩ߻�J������ �'�9���]�o�������$UI_�PANEDATA 1�������  	��}3http:�//1.1.0.�10:3080/�FRH/FCGT�P/FLEXUI�F.HTM?co�nnid=0  �_dummy.h�tm��K�]���)Gpri9�����}������������� ) 7[B�x����v�31p-� 267�Cv�
SYSVA�RS.SV  O�R_PEAKLO�G_OUTPUT�.VR�����  �% ۜ�������  /�$/��H/Z/l/~/ �/�/	/�/�/�/�/�/  ?2??V?=?z?�?s?��?�?�?�?�?
O}  ��)E��E/JO\OnO�O �O�O�?�O;/�O�O_ "_4_F_�Oj_|_c_�_ �_�_�_�_�_�_oo BoTo;oxo_o�o�o!O 3O�o�o,>�o b�O������ �Y��:�!�^�p� W���{���ʏ���Տ �$��H��o�o~��� ����Ɵ؟+����� 2�D�V�h�z���󟰯 ��ԯ�ͯ
��.�@� '�d�K����������� �U�g�%�*�<�N�`� rτ�׿��������� ��&ߍ�J�\�C߀� gߤ߶ߝ��������� "�4��X�?�|��� �����������q� B���f�x��������� ��9�����>P 7t[����� ��(���^p ������a� /$/6/H/Z/l/��/ w/�/�/�/�/�/? ? ?D?+?h?z?a?�?�?�?5G}��?OO0OBOTOfO)�?�O� zO�O�O�O�O�O_xO 5__Y_@_R_�_v_�_ �_�_�_�_o�_1oCo�*ogo�QK�$U�I_POSTYP�E  Q?� 	 so�o��bQUICKME/N  �k�o�o��`RESTORE� 1�Q�  �*default��SINGLE~}PRIM�mmenupage,74,1t ����u��� ,�>�P��t������� ��OuZoя�U��0� B�T�f�x�������� ҟ䟇���,�>�P� ��]�o���󟼯ί� ����(�:�L�^�p� ��%�����ʿܿ� ���ϑ�Z�l�~ϐ� ��E���������߱� 2�D�V�h�z�%�/ߙ� �������
��.�@� ��d�v����O�����������mSCR�E�`?�m�u1sc9pu2�Y�3Y�4Y�5Y�6�Y�7Y�8Y�6�TAT�m� �cQ�j�USER;�@�R�k�s[���3��4��5*��6��7��8��`�NDO_CFG ���k�0�1�`OP�_CRM5  X�5=�`PD������None��b��_INFO �2�Q� �`0%$������ BT7x[� �����/�l��OFFSET 	��i�/��2p�� Y/k/}/�/�/�/�/�/ �/�/E/�/L?C?U?�? y?�?�?�?�?�?;�oMOBO
2OgO��I��WORK �� OVO�O�O/��UFRAM]pV��RTOL_ABRqT_�RENB'_~XGRP 1�-y��aCz  A� }S{Q��{_�_�_�_�_B�V�_�_Z�`UGX�[6[MSK  hJU�6[NQ%�	��%�?�o8U_EV�N&PJd<�f.3ݡ7+
 h[�UEV&P!td�:\event_�user\�o�`C�7�oDO[ FtM�`S�P�a�gspot�weld}!CA6W%7[�zd!zo �o���w2a��� $�Y�����:���^� p��������ʏ܏� g�V���6�H�~�ӟ ������-�؟Q�c��� ���D���h�z��fWf�@3���SA8��!�3� �X�j�E��� ��{�Ŀֿ������ 0�B��f�x�SϜϮπ�����Ͽ����,���$VARS_CO�NFI1 �7+ F�P���3�CMRvcR2�7++i�[ 	\ �B%1:� SC130EFG2 *�߼п��8i�{�2`�S  [�?��P@�Pp�P�N-� �O�� ��;�M�z��u���-�UA�������� B��� �������f�C�� g�R���v��������� <���Q�u��;�GRID�bͪO� �?��}p�>L��@���?� ?,g?�3�3��  @��@F��>��.P������?�IA�D�<�M~�,		��e|WeG�P �x�yH>�ISIONTwMOU�o �����b8�c�rQ FR�:\�\DATA�   �UD�1�LOG�  ��EX���'� B@ �� @"��^/�v/�/��� � n6  �����=!,g�'�5�  =�����!��� -TRAI�N'/�!�"�rd3p�%�(7#KT��{���k (>(9x= 6	x?�?�?�?�?�?�? O OO$O6OHOZOlO�9�IS_GE��n�k�`.P�
wP�.P�B�G$ RE� ��jY��;�LEX�D��� 1-e�V�MPHASE  ��e���>�RT�D_FILTERw 2��k �����_�_�_�_�_�_ �_o#o5o��~_couo �o�o�o�o�o�o�o��	SHIFTME�NU 1�[;
 �<M,%M/c���Ag�w��� �����T�+�=����a�s�����	LIVE/SNA_��%vsfliv�&^ҏ�� S�ETU_���menu����o���R!ub��[9�wMO�m�^�z=�ZD��ɵ�O��<0�@�$�WAITDINE�ND�D1��	�OK�  ��$��?�S�S�&�TIM���~�G���2�ëR�࣪q�����$�RELE=Qӧ��	����_ACT�Ҩ:$��_� �2�%���ӿ8և�RDISt_�T�	�NSP���왴��{�3�z�r�<#�1n:�XVRQ�^��$ZABCz�1��� ,0A�D02ۿ�⑌�VSPT ����$
n�n���N�� �߽�DCSCH��2E0�
A y�-I���@������߹�MPCF_/G 1�<�0�Ð$�6���ÿ��E1pV���A�� �� 18
����Q`� �G۪��Ұ?��J���?�\�?�����?>�����.Il���C�D25D4��0��A@H���*��=���>����{m=���A��Gݛ��g?����Uq��}��ۿ�û�_��.K�������jD4�1�����-q=���>W��������4�� � |�g���>�������Ca~���Տ��:��*����������v��� � )7a����1�57�I�u���P����_CYL�INDcQ�� ��& ,(  *&7##`G�k �����  /p%///[/�/ �/�/��/b/H/�/�/�!??v/W?i?��29���� ��? 4ݗ��?��ON�?AO�ז[AA��SPHERE 2�̻/�O?�O�O�O�O 9?LO'_9_�/]_�O�O �_z_�_�__�_�_F_ X_5o�_Yo@oRo�o�_��o�o�oy�ZZq� ǰ�