��   ��A��*SYST�EM*��V9.4�0341 1/�17/2024 A   ����CCSCB2�_GRP_T � h $CO�MPMATEXP�1 :2F	RI�XU   d$O�FFSEAFGACGEsm;fz�� z_ORG�f � ��P�H F�S_TYTSBF�RAMEe$INIT_TOL��RANGE2_F�f�T�FTR/ATIOe� �_H_LIMU��LFSOFST�_S�mUPS_�����	e� OL_�{UDUMMY2�U�3��4��$$CLASS  �������I��I�VER�SION��  Y5�$�' 3 �I� w���d �� /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"?�4?F?X?j?|?�� �?�  �?�7:׃o�0���@o  'Bd����0@��0 �? x�1EAC�  #E��0�0�09@�Bp�7�?�;VO��FP��