��   ���A��*SYST�EM*��V9.4�0341 1/�17/2024 A   ������CCFR_�LTST_T � x$TP�_PROG �%$DATEJ �$TIMR2SU�F_NUM  w$TlSCHm��CHSoER�Rm  $APPL_TYPR ��ENS�� I�NI_POS� � �FRC�F;IN�MAX�	��DF�F� EMyPq V_LEN,GORI� I .I� �6DUM_R��UL� _FOR�CE_OK�MO�MENTsEND_AVE_F_���OSC_GDW��� _OFST ��/COM9�  $TOT�AL�5 3 o 4/AL� ? x AS ew������ �+=Oas@���1M!: � //&/8/J/\/n/�/ �/�/�/�/�/�/�/?�"?4?F?X?�D9� 8 $� �3 �1P 9(Q4IDX�2�1�X�4�$$C�LASS  ����FQ��'��'�;PVERSION�CX  �Y5�$��dX'���% 	 ���_�_�_�_��s �S��   o��o.o[oRodo�o �o�o�o�o���o �o8J�oOa�� �_��_���oo o!�3�`�W�i����� ��̏ޏ!���8� J���n�a������� ǟٟ����y�F�=� O�|�s�������֯� ���0�B�T�˯Y� v�����埿�ѿ��� �,σ�5�N�Y�k�}� �ϼϳ���#����� :�L���p�cߔߣ��� ����� ��!�{�-� ?�l�c�u������ ��-�� ���D�V��� z�m��߰��߭����� �����RI[� ����%�� �<N`�e��� ������#8/ �A/Z/e/w/�/�/�/ �/�//?"??F?X? �/|?o?�?��?��? �?O/-/�?9OKOxO oO�O�O�O�O�O�O9? _,__P_b_�O�_y_ �?�_�?�_�_�_O%O �_�_^oUogo�o�o�o �o�o�o1_�o$H Zl�oq��_��_ ���o/oD��M� f�q�������ԏˏ�� ;�.��R�d�ۏ�� {����П���� '�9���E�W���{��� ����ï��E�&�8���\�n�寒�������$CCFR_D ����α�'�  ������8�+�=� ��e�wϤϛϭ����� ���"�I�F�X�7�|� ��߲ߥ߳������ ��?�Q��߽ߊ�� ������������]� *�P�/�t�������� ������)���I� [�p��y���� � �$g�HZ9 ~������� 3//D/Se�q/ �/�/�/�/�/�/�/? .?qR?d?C?�?�?? �?�?��?+/�?O)O K/]/�?�?�O�O�O�O �O�O�O�O&_i?6_\_ ;_�_�_�__�_�_�? �_5Oo!o	oUOgO|o �_�o�o�o�o�o�o 0s_TfE�� ����_�?o� +�P�_oqo�}����� ��ŏ����(�:�} ^�p�O������ʟ�� � �7���#�5�W�i� ߟ՟������دϯ� ���2�u�B�h�G��� ����'���ҿ��
�A� �-��a�s���߿�� �ϵ���������<� �`�r�Qߖߨ���� �������K�%�7�\� k�}��߉������� �����4�F���j�|� [�����)������� C�	/Ac�u����� ������ >��NtS��� 3��/M'/9/ !/m�/��/�/�/ �/�/�/$??H?�l? ~?]?�?�?+?�?�?�? / OW/1OCOhOw/�/ �?�O�O�O�O�O
__ _@_R_�?v_�_g_�_ �_5_�_�_OoOOo ;oMooO�O�_�_�o�o �o�o�o�oJ�_ Z�_���?� �o"�Yo3�E�-�yo �o�����͏ߏ� �0�'�T��x���i� ����7��ן��,� c�=�O�t������ ���ׯ����L� ^�������s���ʿA� ���$�[�!�G�Y� {�������Ͻ����� ����)�Vߙ�fߌ� k߰�����K������ .�e�?�Q�9�ϗϬ� �����������<� 3�`��߄���u����� C�����#�8o�I [��������� ��"+Xj�� ����M�� 0/g-/S/e/�� //�/�/�/?�/? *?5?b?�r?�?w?�?��?�?W?�?O$$(+/DOw/UOgO�O�/ �/O�O�O�O�O_._ %_7_d_v_�?�_�_�_ �_�_Y_o�_/<osO 9o_oqo�O�Ooo�o �o�o6An �_~�����c ��1oF�}oW�i�Q� �o�oď�͏��� �'�T�K�x������ ��ҟ�[����,�;� P���a�s�������� ůׯ����:�1�C� p���ş������ܿ� e���3�H��E�k� }ϟ���'��������  ��)�B�M�z߽��� �ߏ�������o���� =�R��c�u�]�ϻ� ��'��������!�3� `�W����ߨ������� ��g�8G�\�� m������� F=O|� �������q/ /?T/�Q/w/�/� �3/)/�/�/�/,?#? 5?N?Y?�?��?�?�? �?�?O{?	O&OI/^O �/oO�OiO�/�/�O3O �O�O	__-_?_l_c_ �_�?�_�_�_�_�_s_  ooDoSOho�Oyo�o �o�O�O+o�o�o %RI[���_� ����}*��Ko `��o]������o�o?� 5�����8�/�A�Z� e������ȟ����� ����2�U�j���{� ��u���ӏ�?��
� �'�9�K�x�o���ߟ ��ҿ������,�� P�_�tϫ��ϗϼ�˯ ݯ7�����(��1�^� U�gߔߦ�����߻�  ���6�)�W�l�� i�������K�A�� ��D�;�M�f�q��� �߮�������
�� !>a�v���� �����K�!3 EW�{����� �//�8/+/\/k �/��/�/�/��C/ �/?4?+?=?j?a?s? �?�?��?�?�?OO �?BO5Oc/xO�/uO�O �O�/�/WOMO__#_ P_G_Y_r_}_�_�?�_ �_�_oo(o�_-oJo mO�o�O�o�o�o�O�O  Wo	"-?Qc ����_����  ��D�7�h�wo���o ����ԏ�o�oO��� @�7�I�v�m������ ����ӟ�*���N� A�o�����������ۏ �c�Y�&��/�\�S� e�~�������ƿ�˿ �"�4ϫ�9�V�y��� ů�ϱϙ�����c� �.�9�K�]�oߜߓ� ����������,�� P�C�t�Ϙ��ϩ�� �����[���L�C� U���y����������  ��$6��ZM{� ���������o e2);h_q� �����/./ @/�E/b/��/��/ �/�/�?o/!?:? E?W?i?{?�?�?�?/ �?O�?&O8O�?\OOO �O�/�O�/�O�O�O�/ ?gO_+_X_O_a_�_ �_�_�_�_O�_o�_ 0oBo�_foYo�O�o�O �o�o�o�O_{oqo> 5Gtk}��� o���(�:�L�� Q�n��o���o��ɏ�� �o$�{�-�F�Q�c� u�������؟���� �2�D���h�[����� �����ӯ����s� %�7�d�[�m������� п�%�����<�N� ſr�eϓ���߯���� �������}�J�A�S� ��w߉ߢ߭������ ���4�F�X���]�z� �ϲ��������	�� 0���9�R�]�o����� ������'���> P��tg����� ���%�1C pgy����� 1/$//H/Z/�~/ q/��/��/�/�/ �/�/V?M?_?�?�? �?�?�?�?)/�?O�? @OROdO�?iO�O�/�O �/�O�O�O?'?<_�O E_^_i_{_�_�_�_�_ �_3Oo&ooJo\o�_ �oso�o�O�o�O�o�o _1_�o=O|s ������=o� 0��T�f����}��o ���o�����)�� ��b�Y�k��������� ş�5��(��L�^� p��u�����ʯ�ۯ �կ!�3�H���Q�j� u�������ؿϿ��?�  �2��V�h�߿��� �Ͽ���������+� =���I�[߈�ߑ߾� �������I�*�<�� `�r��ߖ������ �����#�5߫��n� e�w������������� A�4Xj|�� ��������� -�?�T�]v�� ����/K,/>/ /b/t/��/�/�/� �/�/?(?7I�/ U?g?�?�?�?�?�?�?  OOU/6OHO'OlO~O0�?�O�O�O  