��   ��A��*SYST�EM*��V9.4�0341 1/�17/2024 A   ����CCSCB3�_GRP_T �  � $FS�_TYP3 $�PS_SBFRA�ME3��$J�  $INI�T_TOL^RA�NGE3_F_�uT~FTRAT�IO^c ��P__H_LIMA��L�FSOFSTs_S^JM3_f �_4�$$CL�ASS  �S�����[��[� VERSION��  Yw5�$' 3 �[� 6  � �����D@��  B �� A�����{Cp  T�C;��B�\j�O