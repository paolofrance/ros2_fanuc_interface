��   ��A��*SYST�EM*��V9.4�0341 1/�17/2024 A   ����CCSCB_�GRP_T  � � $COMPMATEXP �9RIX  � 0$INNE�R��P0D_OF�FSETShCsMPAzCOFs�FS_TYCSB�FRAMES  �Y IT_TOL~�RANGE_�� �r�FT_RATIOSh�_H_LIM ��L�FSOFS�T1�
2���4�$$CLAS�S  ����3����(VE�RSION0{<Y5�$'� 3 Q� �<  0 6��S������  a����&Hf��ٸ����� �������  �  BY��� @�  ��� 9!Q%M!C� � a%  �w Bp+'<//�-