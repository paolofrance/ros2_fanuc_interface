��   E�A��*SYST�EM*��V9.4�0341 1/�17/2024 A   ������CC_DI�O_T   4�$D5 YPE�  ?IND�EXGIBIN4�/ MON_DAT�A6  p	�$ENABLF�$BASF   }�_NORMG $LIMIT�|��ERROR����IOCO/ CNTR_CTM}� �$PF�_ENBG 	V�L�PDD_POSRGN%��� LF� CTAPU-a>T�DIS� � FCG��FRQ>/ E�LCPN F} �P$�DTM�ANU �S�ERNO�OPF�L�MODE�S�FTVER���qC_GRP}�d ^$FS_�FORC� ��P>�S_MEA2'%� 1GF#2G0 ��GTSK_CHKZY%O RIc"]!�APP�$PS�_AAML��$�"�	$/!_MI
2�$AS�!!�#�'#�#�!�3  2} ROM_RU2w$J� EST2!�$� �N_NU��$u  3� 
$SB*BS�CNCTOINSv29FS� _NG?$GAGEx� �� CUTFRE�QY#LR*REA�L%� �2MOME�N�T�VC�F2�C��2NC�K1�DT��1DEVIyDS�7 	�3�PATH�0A�3F�NA� )DEXp� �5O �8BUF�7{TD�7COND��;FO_ZD�3CH�G�_@FOS�xAV��7RE�C_TRQ�;CH�_MSp!$LO�C_H�S�Y�FLG�J5�0� � N IU�
@!(UF*����4OSV3EN_yCG"�RTKL��`SSIZtC`SLO�O2!^UD�0iXFLsTY�Z�ZCUR� jW�4@�!�A��Q�S�@1�SMPL.�PEXE����!_�EUR�A��AgXPA@fNE4iT-%0g-(a�AVA?le@Ymd7D�fg�AF���eQ0�EcQwl�gTO�0�H�e7D v�3�e��e�etg�QTP�0I�KS�Q_OP�TCH=IWRR_POaq��ASW�DMM��A@  @ �$�q�EREG_�OFKS�qME�xA1SKS1 Q !�q�RE-   �# �0�r{F�s{Ĺt� M�t ��s$�STD�x��wFA � �x5��w�"��"��/ �q~   �$�pTIN�@��0SUL� �R}_@  $}�@ ys?��O��R�%	 x���0�PJU� ysqFS�4D}
 � �$�0pGF�`qC!$FIL� �@��E�P�A��:�DI\G4�@SCA�8��INTTHRS�_BI�An�SMA9L9�COL����ATE_TI%�P�R�@#��U��!CM�DA	 FSUpEN�V}P $�HRZ_AX��CU3VR�QLB�0����H�����P�NT_MV_AVR�CS5�L��s�C0�v�Cp���ST��x��F�#STO ��F}X�LECTEDC0���Q����FY�����Z���FZ֯w�R�����/ �PO��X $��_I�V����$!0B�"D�?0Z�CCBD�DNQ�CCIw�D?UMMY23G r��DEBU�A\!�PN�"TO��RP"� �c��J�� �;!Ͳ�BUTT`� �@eq��E40N �FS3�a1��T��I%�NEW_UI(ӒV, �U�p~�CCOORD�\GTCH��01P���$%`��~ l ��!�3�PWEIGYHб�2 !�_�q5F��T��WA3a��ƲNTERtaҴ-  �Ů �s���AS0��w$JzASTAа� �q�0�1��*?�2J�3J�W�5�P� ��Ӥ"C�@X��eY��Z��s�CMа�?��X��}�RSL�����Ғ��֢���&��  /�_�~   E0c"0�VROUNDCMV�PERIO˒$Fw1PUU3F2D�'�TM1� �g�_D<IcGAMMc1Jb��TRX�eK��K��K��CL��&On00ADJ�GA�CUPDC�R6���E�S��QREX���FR_� @W��&�#�u2�DL_R��T�Q�MXp�3x�0���#�� ���"���� �����������������VL ~�6,
��UK��tD,
`�P5A8@W`
X�A� �6 �y"��gVIBڶ�OV�
DEH�栐�p@�)�@��>�)� ��RTn��MN1HS;vMN2mUFRA���9x�zA�`A[���OR�`(��AL%�!��CJ��`�&�6S�8B�I˅L .$M˂P30?#�a =$�`�˂��$HCcB$�GV��GV��GV��JDO��q��%S.�#$R&�E��r4�#q�U�AP=�DA9�$�3$V�P��b�1Lj ��(PIL�� U��!��3��2�@Wb�5��OA�?���!�V07�!�5OBODA@��Y�MR9G7A	�4��453��E([��p�;�uCNPRG�OVJ��5�P�_T�W@�BG?�E�M�NVfcD��DWT��sk�TRL_SK�I~�JyqIcN��G�WJ��eRPENA�BZ�j�j#5 ?� A$SB�� 0cɓ��3`��1b >�,h�1bXQh4�/�&��B_KQ��S����%ALARMSERua� UTOT+TFRZGCHKE%�����F2�IbS�DbP�E2pbP��J�Z� �U�B2�K2p�MbQMU�VFIXF�"�RF����(PI�tX��� DON��I��SyFg�@_DF165BF2Co�Zɐ���DR��P���C3Q��E ��X���Z�j� �e�B�3�K3�M��MU�cD�IA�0�Fr_��R�
v�Uv�S�CGA�P�P��rPyjAPt ���`v�au�ev�cC$���0$��VU'"z�UD��S_HA�aU �u�t�DGEZ  �@�B�p�K��%�E55u,�_�53�l�4!	ԃ���m��q0��_FSIW4! W� >�X��R_���pHK�_CHC9K�1;�INSA0���0PReO0ˊH�NT���̉�Qt6�������d��� ������$����8����4F�Q�Q� ;�� �SIOy�E�  Y5���}C�BSV 3F��~�� � � )�������Ú@�Ù	������F@� �Ր��8�  Q�o�I�W�i�@{���������Q�dQ�
Ӡh���ݯ�� ,�N��F�M�L�F�X� r���ˢD�v���¿ؿ ���� �.�\�
�d� NϤϚ���v��Ϻ��� ������N�`�z�<� �߀������ߨ���� B�8�f���X��� n���,����>��-��?�0�	UD1:� 678  A�fsdt1 789012345h�xw�����  )o�0g������.����N�R�'G���� l�+�H�` 71�u����c�O����� ��LCU�y ������/��6/H/  u�DMM� d���K,A  []�/�/�/�/S+�`�OR 3	g+ Q�u�nAZ����B?��o�4-2S4D 
g-!n�o?z7���?��?���(� ?��#B���0���)**�*�?�?�1�?O�/C���ONFIG �F����M�2�.D��.Oϡ��D  �z�  D�@�E��!�R��@���Co  CuC��A��uBDDk�/�2uCN @C�.� 3<,`��_�/-_Z�ͣ�=���A�1 �-2/u_�_�_֟�_�_ �_o�_2ooVoAozo�@�j�c�o �o�o�o�o�o
. @Ryro�r���@����)�[#Iz�� 3g) AQ�Z�`�fQ,���0��oPB�1��nQ�C��@����=#׽
��Nnk(��K������U@��=e˅=D��ׅ���;����8I�y���It$ ��$,�kE��I��7�Fۀ3C�jR�_��_w�n�����+�{�̫�.��������$敕Ǖ(4�$�ӕ����>�E=���B<~w����8E�y�;�j�'�ǂ��7�>'��C���?�0S��z�BHY��1�0>���fQ@h�_���.���Ȣ@.��F��3Fs�"ǔ�E�ȯ+�C���C�B��B�����1bjQA�1�1|�Bp�3�B����1ۡ@۠@4h��0@�@@�k��! ���"iG��o�o�e�ҿ ɿۿ�w���C�fR�0C���?Z�O��0C�<�?�33k�}��:�o�ϥ�� ��������k��͘w�@�n�?Lm�]!S�C�<8< ��ќW�X�W�V�B����2��@�������CX������ �1��ߢߤޓB�� ���߄�
��.���L� n�$����K���e�� ��2���A� ��@����%��C�<@��P�L8�g^]o���|� x
l�G����-@�Y ���0h���v]!�_FCCOORD� 3g+2 `! _�>/��I/ �/p/2/�/V/x/�/ �/�/�/�/$?
?�/i? ?>?�?R?�?v?�?�? �?O�?ODO*OO�O <O^O�OrO�O�O�O
_ �O=_�O"_d_J_8_�_ \_~_�_�_o�_�_*o �_]ooBo�ojoXo�o |o�o�o�o#�o�oJ }0b��x� ����C���j� ,���P���ď����	� ��ޏ0��c��8��� L���p����ʟ��)� ܟ��P����6�X��� l�ݯ��¯��دI� ���p�2���V�x�ʿ �������$�
���i� �>ϐ�R���vϘ��� ������D�*�߉� <�^߰�r��ߖ߸�
� ��=���"�d�J�8�� \�~���������*� ��]��B���j�X��� |�������#����J }0b��x� ���C�j ,�P����	/ ��0/�c//8/�/ L/�/p/�/�/�/�/)? �/�/P??�?6?X?�? l?�?�?�?O�?�?IO��?OpO�C�$CC�_FSIW �����A��  �F�H�A�L�O�OT