��   F�A��*SYST�EM*��V9.4�0341 1/�17/2024 A   ������CCHG_�LIM_T  � �
$COM�MENT �$CTRL_STATE  M�IO_TYPX
I�DXXUFRAM�E_NUMxTO�OL�INSID~WMARGINX �$UPP_XY�Z4   �$LOW�4/C�FG8� a�$KNOB_MO�UGZ �SE�L�EF�GRIP_wENBOPE� {)CLOSW �)LEVER�L�V_DIR_PY�XBTN_OUT�YeYuONE�_HANDXAV�G_F�� ROT�_^TRNS� T�R �b�uSFD�OD�  �$ORG_PTH�_RES�TOUCH�OC�*��$JNT4MR�G�3$,$�G+C"2a3�U"l(�SP�8u#�)�WPR�*�)�DC���#$R�EC_METHO��'b �$e�$uT�EACH_PAT>#MULTI7�!|�&CUSTO��GEN_TP_PRO= )T�*�� �e=�� ]1DEV��5���_AR� 3  
�K9_2 �K_S0�n�1ENC�SB~�2,$�0_RIGH��/!HDL_MAS�BCV1�A�2�VA�5EG�5E+L=JML+G�1F_�1 �7�FF_VAL�ID_M�MAX�_RUN� + � GAIN��G� �3!�� J(k!�F� SNG�L�R;"��B� P���X�22T�!�0_AR�3�!�PT]1C��CUR_F5PTS�M�@wX�APUSH_F�C�@�Y�U�T�Uħ3;T3S��'$�!�YJ1_R�V�@�j5�[SIMPLE-QXOF�F<a�E3SH� M1OK�^�.RO�RSV Nt� �2sbREA@ܻ�cSTR|a?>�0DEBUG� ���DATA8$ S�6�@ ^�@ �esP�oT�lb.*� rQ3!wrl lc�02�S PRSW�NE��REBO�2�I�T�]dNON_R�ST�FSA/bITgnsORCW ."�r��C."MEAN�zH�DGD_ACTI�VWSAFEM1
��tO�u�r�@�$0�`�X�P PS�T�bNEqp�4 �S�S�xf�S_W�P."EX�{ -�h�,$��@�`�V] ��3!�!��l ���T�� d��d��-���X����SMAL�A���@OCVR���+��FO=���@l H�1G�U�5�G�BE���vAF���wESCAPE��TOP�f$CL�AL�aAlTDDS1BrQ�!TCg � �e�%rQ�)rS�Wꕿ)  Yu�"*z�w���������rQ.XM3?V?uE�gSUBS0GtN�O_M�Ė�DBp=!ߦȦ�WAIXt��jP�A��b�'8�NiT`r�qbT_ϓ:Y�C�DOW3Sm�1N�v�3�FC���1�B�e�1T @�gtfV���jV�2/ MQ0� 6T��P�9Vmd ]l`@0yA`�.���!T�dTL_OR84 �E�AMOMW�2����GRV_OF C2���!�2��`F�ÇRSL��LQu!�F!I�q�$ud��f�����GRP>8 A
T4%$Dqp��II2O�R8��1DI��3aAPW�3�5VE)@�E�7jՄj�OCIiTSjVR@0MD�' �jѧܠQ2v}�@���Sp���B�bS��\ 9$PA�US����G�AB�WҔDAP5 	U�oq���PW� W0M��@z�FIb����U���ERR �f���BdW���RETRY%�,Q�� �������T`HtC�%AqpR�A3�O�1�3�BՔ�1�\��]�b���W\Tpb0��u�rLO�b]�?���LOO����"2�������+�������EN�5d��Y�E���P]�Ua�U`RT�\Ǖ3�ONLSP� �OFFG�BLIN �1c�Ė��� w�B K�7UaALAR���Q�)�q�� Ua�КҦkX�)'�bx��rn�Ǎd�eP(�Y�W���ӑh=���O*�ID1`�H��h�,OPER����I���P�C�_~@	$WIR`p��sPC��"� ���9!CHAR�:�VOOLTAO(�CҖ�RI*�O�;�O�a�Lr0�`0���?CONNECL��6OT�`�����-"0Ґ���A�&NE{�S �3꒼aM��"6��� ���6.�� �S9,d3PA��"T��i6�1w7�aIN�p!�4�0�4] �7] �3�daj3!��PATH���!~b�cTt�`X��8�bs��;Js�@��CsPZ!EH�I~ �,a�zʼrV��Ê�aD�1�G�1�H3�K4�K5�A �$�̑SS6����4�A5�Y5� Y�@�PoSION�H���Y5�$�b� �XY��A<Y) �AP_b_I_�_h[���_+B�hV�V�P�_ΧU �_hU@��5��PF< o<�b�`0oc4aCH'  A`Ta@�_gm�R)
��!�_01h�_�n�Q�A?�
d?
 P �o�S�]BQ`/�E;� �e�a��`u�o �o�o�o"4FX j|������ �[��0�B�T�f�x� ��������ҏ���� �,�>�P�b�t���hZV�PBζT��P��T�����?�3�@ ��  �X�P�Qɐ�UA�*�<��`W��ȑ���UaĽQA��M�L��`=����L�BM�=L���?�p�P�� B aɐPb��ء@�դb u0  Ь�.��  d\a>�a��=?��<#�
H�Yd �b	e5ਦ��2�_[� m��������ǿٿ� ��D�!�3�E�W�i�{���ϟϱ���hX
 y_hR�����1�,� >�P�y�t߆ߘ����A"T
1 /Y�a� �������.ﭙ�_�[ P�ﱛ�����hZ�����6�H��� Q�~�u����������� ����2D��F jq������ �� �9K2o� �������/ #/5/|�k/}/�/�/��/�/�/�/�/?��MkTP(S/\'����O0�ǐ�W?�T L?�?�?�?�ِ?�?O�O?GRP 3�/[2 ��� %s	M�o}O 	'0��qL0?�
`\`ܢ N)�hX�AUOgI�A _�OZ�O�O�O�O�O03w__�@�Z8_J_\_n_�_04o�_�@�#j�_�_�_�_o05 �o6o�@�jXojo|o�o�o06'�o�@Cz�o0�o007�V��@�zx����08G���@c���,�>�P�09׏v��@� ������Ώ��1󠅟����(�:�L�^�p�1 sO�����O��ϟ�� u�_%���+_M�_�q� ��u��_�����_ݯ� ��u�#oE���Kom� �����u��oտ���o ���!�3�u�Ceϧ� k�ϟϱ���u���� ����/�A�S�u�c� �ߧ����߿�����u� �六�=�O�a�s��J2����@"����������2�5�G�;� ]�o����������G� ˯����#�3�U G�[�}����ÿ �G��1C� S�uG�{ϝ��� ���/G��-/?/Q/ c/�sߕ/G�߽/�/ �/�/��%?G�+�M? _?q?�?���?G�� �?�?OO�J3#�EO�'P�KhOzO�O�O�O3 ���O�A���O_!_3_ �KCe_�Ak�_�_�_ �_�K��_�A�o/o AoSo�Kc�o�A��o �o�o�o�K��A/ =Oas�K�/��A �/�����K?5� �A;?]�o������K�? ŏ�A�?����#��K 3OU��A[O}���������4�O�Ǡb���,�>�P�4S_u���{_ ������ӯU��_��� o-�?�Q�c�U�so�� ���o��Ͽ��U� %χ�+M�_�qσ�U� ��χ�������� U�#�E߇�K�m�ߑ� ��U����߇�ۏ��� !�3�U�C�ek��� �����U�ӟ��� �/�A�S�5
5c����g ���������$�CCSHG_CF�G ���>�Y���mU����a�
�������B� �������� a����������' $��f����������/1/C/U/q	� A ��	Z/E	1?234567�����%90�#�/�!�/�	?���!�+,?  !�-\;LT?f? x?�?�?�?�?�?�/�/��O4OFOXOjO |O�OX�O/�O�O_��O�OC_U_g_�� �?�1�_�_�_�_�_�3