��   ��A��*SYST�EM*��V9.4�0341 1/�17/2024 A 	  ����DRYRUN�_T  4 �$'ENB � $NUM_P�ORTA ESU�@$STATE� P TCOL_���PMPMCmGRP_MASKZ}E� OTIONN�LOG_INFO�NiAVcFLTR_EMPTYd $PROD__ �L �ESTOP_�DSBLAPOW�_RECOVAO{PR�SAW_� �G %$IN�IT	RESUM�E_TYPEND�IST_DIFF>A $ORN41p� d =R�4&�J_  4 �$(F3IDXX��_ICIg�MIX_BG-<y
_NAMc gMODc_USd~�IFY_TI�� �MKR-�  $LIN�c   "_S�IZc�� �. �h $USE_FLC 3!�:&iF*SIMA7#Q�C#QBn'SCAN��AX�+IN�*I���_COUNrR�O( ��!_TMR�_VA�g# h>�ia �'` ����1�+WAR��$�H�!�#Nf3CH�PE�$,O�!PR�'Ioq7�iOqfOoAT�H- P $ENABL+��0BTf�$$�CLASS  O���A��5��=5�0VERS�G�  Y�@'/ E5�������-@]F!@AbE��%A�O���O�O����3EI;2>K �O_ /_A_S_e_w_�_�_�_ �_�_�_�_oo+o�O�)W?"HI@ ��lj@|o�o�i��� � 2>I  4%:o�o��_AoA�o�oAS 2w�h���� �i
B���j�I��{��{�c$"+ �ktK-@b����bA��X_A A-@vNڏ����"� 4�F�X�j�|������� ��bFoAǁoA���
� �.�@�R�d�v����� ����ЯDZM���@�7 2�lǏ1� C�U�g�y��������� ӿ���	�Ɯ#�<�N� `�rτϖϨϺ����� �����8�J�\�n� �ߒߤ߶��������� �"�-�F�X�j�|�� ������������� )�;�T�f�x������� ��������,7� Pbt����� ��(:E^ p�������  //$/6/ASl/~/ �/�/�/�/�/�/�/?  ?2?D?Ch�4�0��{? @