��   ?3�A��*SYST�EM*��V9.4�0341 1/�17/2024 A   ����MN_MCR�_TABLE �  � $MA�CRO_NAME� %$PRO�G@EPT_IN�DEX  $OPEN_IDa�ASSIGN_T�YPD  qk$MON_NO}�PREV_SUB�y a $USER�_WORK���_�L� MS�*RT�N  4&S�OP_T  �� $�EMG�O��RESE�T�MOT|�H�OLl��12��STAR PD�I8G9GAGBzGC�TPDS��REL�&U�s �� �EST�x��SFSP�C���C�C�NB��S)*$8�*$3%) ''5%)6�%)7%)S�PNS�TRz�"D�  ��$$CLr   O����!������ VERSIO�N�(  �Y5�:LDU�IMT  ���� ����$MAX�DRI� ��5
��$.1 �%� � d%
�Vacuum O�ff����K0ACU?UM_OFFa?��K	���!��q0=	M5n  1�?k6!	u5� �?�7.�6�0��4Relax �hand�?i8 $)OOO �"�3�#q0_OpenC2QO�2O�OVO�3 qDClose}O�O�O_bI�GH�O�Oo__�3oFh_�_d_�_�[ �3�5�_o�_=o�_�_ so"o�oFoXo�o�o�o �o�o9�oIo 0�T�x��� �5���k����>� P���׏������1� ��U���P���L��� p��������ʟܟ� c����6�H���l�ͯ 󯢯��)�دM���� ��2�����h�z�￞� �¿Կ!�[�F��.� @ϵ�d��ψϚ���!� ��E����{�*ߟ�N� `ߚ��ߖ�����A� ��Q�w�&�8��\��� �������=����� s�"���F�X������� ����9��] X�T�x��� #��k�> P�t����1/ �U///�/:/�/�/ p/�/�/�/?�/�/)? c?N?�?6?H?�?l?�? �?�?�?)O�?MO�?O �O2O�OVOhO�O�O�O _�O�OI_�OY__._ @_�_d_�_�_�_o�_ oEo�_o{o*o�oNo `o�o�o�o�o�oA �oe&`�\� ����+���&� s�"���F�X�͏|�ݏ ���ď9��]��� ��B���ɟx������� #�ҟ�1�k�V���>� P�ůt�鯘����1� �U�����:���^� p��������ʿܿQ�  �aχ�6�HϽ�l��� �Ϣ�����M���� ��2ߧ�V�hߵ����� �����I���m��.� h��d�������� 3�����.�{�*���N� `�����������A ��e&�J�� ���+��9 s^�FX�|� ���9/�]/// �/B/�/f/x/�/�/�/ #?�/�/Y??i?�?>? P?�?t?�?�?�?O�? OUOOO�O:O�O^O pO�O�O�O_�O�OQ_  _u_$_6_p_�_l_�_ �_�_o�_;o�_�_6o �o2o�oVoho�o�o�o �o�oI�om. �R������ 3���A�{�f���N� `�Տ���������A� ��e��&���J���n� �������+�ڟ�a� �q���F�X�ͯ|�� ����'�֯$�]��� ��B���f�x�ſ��� #�ҿ�Y��}�,�>� x���t��ϘϪ�����C���� %
Se�nd Event�U�5�SENDEgVNT��3�	�i�� %	}�Datya�ߘ�DATA��ڿڒ��%}�Sy�sVar��SY�SVY�ڔ1�%�Get��Z�GE�T��%R�equest M�enu����REQOMENU!��ۖ�� ?߀�;ߤ�_������ ������F��j +�O���� �0��fxc� K]������ >/)/b//#/�/G/�/ k/}/�/?�/(?�/�/ ^??�?�?C?}?�?y? �?�?�?$O�?!OZO	O O�O?O�OcOuO�O�O �O _�O�OV__z_)_ ;_u_�_�_�_�_�_o �_@o�_o;o�o7o�o [omo�o�o�o N�or!3�W� �����8��� n���k���S�e�ڏ�� ��������F�1�j�� +���O�ğs������ ��0�ߟ�f������ K���ү��������,� ۯ)�b��#���G��� k�}����(�׿� ^�ς�1�C�}��ϵ� �ϝϯ�$���H���	��Cߐ�?ߴ�c�u��$�MACRO_MA�X:�������Ж��SOP�ENBL �����՗�r�r��A���PDIMS�K����Y�S�Uc�u�TPDSB�EX  -�q�U����n����