��   u�A��*SYST�EM*��V9.4�0341 1/�17/2024 A   ����CCSCBG�_GRP_T �  $SE�RIES_TYP�E  $PS�_PRM_UPD�A��I OTE$�MODEL_NA�ME :An O�tNSWEIGH�T $DIVC�ONST_FF z�T�SBFRq�  $RA'NGE� ��� ����P_H_LI�M��L�FSO�F� S��M_I�NI�DOU� R{EQ�DIGI��+��$$CLA�SS  ����P��u��uEV�ERSIONM�  Y5��$' 3 nu��F � 
W ������� ���� B  y ��C�  %�Bp��!/N/  