��   ��A��*SYST�EM*��V9.4�0341 1/�17/2024 A   ����CCPTP_�CFG_T  �h j$DAT�A_PATH �!$OUTPU�T>5$PART�_NAMEC $�EDGE\!$C�LR_VDB_BUF  $x�_SIZ 9V�ER�DEV_I�D�H �VIS_�RES���P_D�T�POS_OF�S_ENB�TA�R_D� �CHK�_f �MANUA�L_BAK�EB?UG_MOD` X_FC_PN��.�5CUV8S�EG8LAP)TPP_� )X)fH�f�A�� L�WAIT_TM �$ABV_PT�H���RETRsEA� �CNS� ��JUMP_LE�N_�$CURQV)u�T'T)�MAs'ABOV�E_��$TO�L_WPR_CH�gn!q EXP%S�Ac A�ERR_H���-����(��_PROgE N�ON� OP�CF%_b R� 4Rf 4�DI� 4LI�D?EACT_F�<5�5XID6�6J8 t9LOC6" ȶ5�P��AN�0�$XD!A���4�_C6CO!�5F�IR �0W�SQ�0Xwn#fj'�E`WO!��$N_� 9L�!�ACHII��L� �DYN_CO SW�JH�Xp�!�: �ALL�
�EP�TW@�
�D%�F�NU��C��A8.� VBASFW@&�XY-Z,WSW@�I��0@0-Z�SPUS X@ViI2U�~VX2oGAINVXYRQ��F�P�Y�P�5}0R6�MI EC�.��Xk;S2CMDp� ~�KANG1Bj	2Bf�LOa�!ec]a�� S% L`_C �  ~bga�b� &:1 L� �3]3�6�TO�T��c��AV�G!�$3�FINI zA�G�yUze@�F�6�Q�3��dU�Dt� �`
BsENT��`7b�y�b�3e�v�f� �k�q�`~bST��  ? 
��4�$s ASS  ���
����Z��Z�p� SI�ON� ? Y5�$'2 �(�Z�!FR:�\) \����5UGD1:]������Ĵ���!��ޏ���A ��3���
���N���u0  �(� �d��(���3�  �@@B�G�?���BHJ�Y��  >�i�`��f���`�Ȃ�*�����Ɵ���B�џ��	�h�`�A&��Dz������֛��?e�H�u�t�H�M�Fl�,$�\���2��!��������ů ׯ������1�C�U��9�:�`G�V�����
�˿������� (�:�L��pςϔϫ��1234567890����� ������ ��$�6�H� Z�l�~ߐߢ�