��   #��A��*SYST�EM*��V9.4�0341 1/�17/2024 A   ������DMR_S�HFERR_T �  $O�FFSET  � 	4/GR�P: $�MA��R_DON�E  $OT�_MINUSJ � 	sPLzdC�OUNJ$REF,j�PO{���I$BCKLSH�_SIG�EA�CHMSTj�SsPC�
�MOVn �~ADAPT_I�NERJ FR�ICCOL_Pz,MGRAV��� HISID�SPk�HIFT�_7 O �N\m�MCH� S��ARM_PARA�O dcANG�o y2�CLD�E7�CALIB�Dn$GEA�R�2(��� RING��<�$]_d�REL�3� 1  	��P CLo: �� �AX{  �$PS_�TI����TIME ��J� _CMD,��"FB�VS �&�CL_OV�� F�RMZ�$DED�X�$NA� %��CURL�W����TCK5�wFMSV�M_LIF	��`;8G:w$�A9_0M:_��=�93x6W� |�"�PCCOM���FB� M�0�M7AL_�ECIr�PL!�"DTYk�R_�"�5L#�1EN�DD��o1� �5M�P PL|� W �  $�STAL#TRQ_�M��0KN}FSD� �HY�J� |GI�JeI�JI�E#3AnC�uB�A�4�$�A{SS> ���	Q������@VER�SI� W  Y5�$S� 1'X ���� 	 ���n_Y_�_}U{�5��9N2��3�M�[|��}'�!��X_�_�|W5  9N� 
�3 �? |� �\�S 2P�T.g,e|YQToBl���r��S�J�s�Ǿ���o�p�� Ao�o�_gl�o�o�o�q�� *< ̟fp�$7w�g �@BNpSp �@
Yu�o�su����t���W����Px n���dw�����=L3���.�?�/���@�O�t��������� Ώ�����(�:�� 	Ue�s�]���T  2�ğ֟������0�B�T�f��R ��������Ưد��� � �2�D�V�h�z��� ����¿Կ���
�� .�@�R�d�vψϚϬ� ����������*�<� N�`�r߄ߖߨߺ��� ������&�8�J�\� n������<��� ������&�8�J�\�n������|(u��q ������2/h S�w�����v
�$&4 1D\���N��K��ZwK�mbL��I�L�:L��P�A�*�B���BOZ��>ʺ�?)��>\�z�B� � �����lB��qs���y��o��>�=�GV�fHE�\Cm�?���@
n?��~D�/��>xFgJ�N<zRTU�UL���g/��/v/�/T�(U'���!�(�/V�� � � L�h���B�&��;ܾ��7��o@>=�����B�����������oI>=N�-�=���Rj��@�-X>��Q�����=���R�� �]�%PAYLOA-�??h�3���BB���_�X��i�2�oCu>=���*?��B����B��	���o]>=���-<9C�+�@�n=����\8�<(� ��?�?bO�?3U"��KB�p�r����n�Q>��B�Y�[�D���f�o��>=��-;
�(k��l'?��3<���ݿ�ϙ���x?JC	rRO#_vN ���/`_ K_�_o_�_�_\�_�_ 6_H_o�_=o(oMoso �_�_�o�_^o�o�o �o'9�o]�o�o� �����R#� v�Y��}�h����� ���<����
�C� .�g�y�̏�����ӟ N�П	���-�?���c� ��ȟ�������ͯ� F�X�)�|�ޯ_�J��� n������ݿ0�B�� ���I�4�m��ҿ�� �����T������3� �Ϙ�i߼�ߟߊ��� ������L��p߂�S� ��P��t������ 6�H����=�(�M�s� �������^����� ��'9��]����� �����R# v�Y�}h����|H����
/ ��$PLC�L_GRP 1����;!?� pzB0�?�  T*l>�?m��T)��/� �/�/�/�/�/�/�/+?�?O?:?s?Z?T.�? 