��   v��A��*SYST�EM*��V9.4�0341 1/�17/2024 A   ����UI_CON�FIG_T  �x L$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�73�ODE�
4�CFOCA �5VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j �Ơ!BG�#�!hIN=SR$IO}7�PM�X_PKT�?$IHELP�� ME�#BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�<S�TYf2$Iv!_8Gv!k FKE�F�HTML�_N;AM�#DIMC4:1>]ABRIGH83s oDJ7CH92%!FEL0T_DEVICg1�&USTO_@ � t @A�R$@PIDD�BC��D*PAG� ?xhA�B�ISCREu�EF���GN�@�$FLAG�@�4&�1  h �	$PWD_ACGCES� MA�8��hS:1�%)$L�ABE� $T�z jHP�3�R�	>4SUSRVI 1  < `�R*��R��QPRI��m� t1�PTRIP��"m�$$CLA~SP ���a���R��R `\ SI��	g  �Y5�$'2 �I�S��R	 /,��?���aa1`jbed`a����� ?�  cd�o��
 ��a�o�o �o%7 �o\ n����E�� ��"�4��X�j�|� ������ďS����� �0�B�яf�x����� ����O������,� >�P�ߟt��������� ί]����(�:�L� ۯp���������ʿܿ�a`TPTX����l��� s� �鶄�$/s�oftpart/�genlink?�help=/md�/tpmenu.dg޿xϊϜϮ�g�9&C�U�pwdd��� ��1�f�U�g�yߋ� �߯�>�������	�� -����c�u����,�����a�`���b�� ($R����`��6�!�Z���a�da��c���c��~�N��k
��da��a�a�J�  ��J�	.H������跦�q�`���`  ����H Gp ���K#J�Ffbc �:c�B 1z�+fR� \��_}�� REG V�ED?���wh�olemod.h�tm�	singl��doub�tripbrows3b� i{�W������"/����dev.s�lo/� 1r,	t�/A�// K/�/�/?�/5?G?Y?8k?}?�?� ��? �?�?�?OO+O=OOOaOjE @�?�O�OpO �O�O�O�F�	�?�?_ /_A_S_e_w_�_�_�_ �_�_�_�_oo+o=o Ooao/'yoso�o�o�o �o�o�o1CU gy������ �? �2�D�V�h�z��� �����O���Ǐُ .�@��O	_������� ��П˟ݟ���%� 7�`�[�m�������� �oկϯ���!�3�E� W�i�{�������ÿտ �����/�A��|� �Ϡϲ���������� ��B�T�#�5ߊߜ� S�e�K��������,� '�9�K�t�o���� ����������߯1� +�Y�k�}��������� ������1CU gy��k����  2DVhzu� ��������� �@/;/M/_/�/�/�/ �/�/�/�/�/??%? 7?`?[?m?;��?�?�? �?�?�?�?O!O3OEO WOiO{O�O�O�O�O�O �O�O�4_F_X_j_|_ �_�_�_�_�_��_o��_�_BoTobj�$U�I_TOPMEN�U 1-`�a�R 
d��aQ)*def�ault_ ]�*level0 =*[	 �o�0��o�o�o	rtpi�o[23]�8tpst[1=xY��o�o�=h58�e01_l.pn�g��6menu15�y�p�q13�z�r��z�t4�{��q�� ?�f�x���������R T������1�C�҄�prim=�qp�age,1422,1J���������˟ ֏���%�7�I�ؖ�^�class,5R���������ϯڔf�13֯��0�hB�T�ۓ^�53p�@������ƿؿۓ^�8��%�7�I�[�ڟ�ϑϣϵ�����Y �`�a�o��mΙq�;�Y�CvtyN}6HqOmf[0PN�	�Пc[164=w��5�9=x�q)�o���x2 ��}Q����w�{�� O������� ��$� o�H�Z�l�~�����1� �������� ��e�22gy���> p���	-�� ��n����e�w�1���//*/</���^�ainedi�	�s/�/�/�/�/���config=s�ingle&^�wintpj��/??�*?<?����r?!ٙ�gl[�ڔ�?vߔ0�8���1���?O�82 ��&O�?EOoO�z��z�4s�x�O�O �x��ON�'_9_K_]_ o_�_���_�_�_�_�_ �_o�_5oGoYoko}o�o�$;�$doub��%oc�13~�&d�ual�i38��,!4�o�o�o9�o�n �o�ax��#o� ������>�P� b�t�����O�a�bڏ ����"�-�F�X�j�|������J]?ҟ�@/�UE��O���s��:�_���G�u����� n�l��O�O�,�R�@�6G�u7��� ��ÿտ�2���/� A�S�e����ϛϭϿ�P�������"�1� /�A�S�e�w߂ϛ߭� �������߄��+�=� O�a�s�������� ��������6
�?��Q�c�u����$��74������������C����6�	TPTX�[20�=aAY24 G,���BY1�8� �����8tHt��`aA��=��tvB�H4���@2p-0��11pi�S:�$treeview�#��f3��Q}381,26�o//A/S/�w/ �/�/�/�/�/`/�/?�?+?=?O?�o���5 �o%���?�?�?�/O O)O;OMO_Oj?|?"	2�?"2-��O�O�OxO��1�?�E��H_Z_�l_ �6�O��edit�a _2_�_�_�_ ������_�C�_Qoco uo$vo�o핪o#�o {�o�o1CU z�os����� �
��y�3�Z�l�~� �������?؏����  �2���V�h�z����� ��?����
��.� @�ϟd�v��������� M������*�<�˯ N�r���������̿[� ���&�8�J�ٿn� �ϒϤ϶���wo�o�� �o"߉'�E�W�i�{� �ߟ߱���1������ �/�A�S�e�w�9��� ����������e�>� P�b�t�����'����� ������:L^ p���5���  $�HZl~ ��1����/  /2/�V/h/z/�/�/ �/?/�/�/�/
??.? ����d?߈?�ߍ�? �?�?�?�?OO)O�? 5O_OqO�O�O�O�O�O �O��_&_8_J_\_n_ �_�/�_�_�_�_�_�_ �_"o4oFoXojo|oo �o�o�o�o�o�o�o 0BTfx�� ������,�>� P�b�t�����'���Ώ �������:�L�^� p�����C?U?ʟy?� UO�O�#�5�G�Y�k� ~�������ůׯ��� ��1�C�_z����� ��¿Կ��
��.� @�R�d��ϚϬϾ� ����q���*�<�N� `���rߖߨߺ����� ����&�8�J�\�n� �ߒ���������{� ��"�4�F�X�j�|�� �����������������*defaul�t؞*level8a���Y�w��! tpst�[1]�	�y�tpio[23���u�d�,>�menu7_l�.pngA^1	3cp5x]�[4�u6cp��� 	//-/?/��c/u/�/ �/�/�/L/�/�/??�)?;?M?�"pri�m=^page,74,1R?�?�?�?�?�?�"f6class,13�?OO 0OBOTO�?�25ZO�O �O�O�O�O�#�<~O�_$_6_H_Z_]?o218v?�_�_�_�_�_�O�26�_o-o?oQoco�B�$UI_US�ERVIEW 1�����R? 
��jo��o�o=m�o�o	 -?�ocu��� N������o$� 6�H����������ˏ n����%�7�I�� m��������`�ԟ �X�!�3�E�W�i�� ������ïկx���� �/�A����`�r�� ����ѿ���Ϫ�+� =�O�a�s�ϗϩϻ� ���ϊ�����߂�K� ]�o߁ߓ�6߷����� ������5�G�Y�k� }�(ߊ��� ����� ��1���U�g�y��� ��@���������	�� ��(:��^��� ��r�); �_q���R� ��J/%/7/I/[/ �/�/�/�/�/�/|/ �/?!?3?E?�R?d? v?�/�?�?�?�?�?�? O/OAOSOeOO�O�O �O�O�O|?�O�O_tO &_O_a_s_�_�_:_�_ �_�_�_o�_'o9oKo ]oooh